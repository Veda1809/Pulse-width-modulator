magic
tech sky130A
magscale 1 2
timestamp 1700890851
<< obsli1 >>
rect 1104 2159 12788 13617
<< obsm1 >>
rect 14 1980 13602 13864
<< metal2 >>
rect 13542 15266 13598 16066
rect 18 0 74 800
<< obsm2 >>
rect 20 15210 13486 15266
rect 20 856 13596 15210
rect 130 711 13596 856
<< metal3 >>
rect 0 14968 800 15088
rect 13122 688 13922 808
<< obsm3 >>
rect 880 14888 13122 15061
rect 800 888 13122 14888
rect 800 715 13042 888
<< metal4 >>
rect 2404 2128 2724 13648
rect 3064 2128 3384 13648
rect 5325 2128 5645 13648
rect 5985 2128 6305 13648
rect 8246 2128 8566 13648
rect 8906 2128 9226 13648
rect 11167 2128 11487 13648
rect 11827 2128 12147 13648
<< metal5 >>
rect 1056 12672 12836 12992
rect 1056 12012 12836 12332
rect 1056 9816 12836 10136
rect 1056 9156 12836 9476
rect 1056 6960 12836 7280
rect 1056 6300 12836 6620
rect 1056 4104 12836 4424
rect 1056 3444 12836 3764
<< labels >>
rlabel metal2 s 18 0 74 800 6 PWM_OUT
port 1 nsew signal output
rlabel metal4 s 3064 2128 3384 13648 6 VGND
port 2 nsew ground bidirectional
rlabel metal4 s 5985 2128 6305 13648 6 VGND
port 2 nsew ground bidirectional
rlabel metal4 s 8906 2128 9226 13648 6 VGND
port 2 nsew ground bidirectional
rlabel metal4 s 11827 2128 12147 13648 6 VGND
port 2 nsew ground bidirectional
rlabel metal5 s 1056 4104 12836 4424 6 VGND
port 2 nsew ground bidirectional
rlabel metal5 s 1056 6960 12836 7280 6 VGND
port 2 nsew ground bidirectional
rlabel metal5 s 1056 9816 12836 10136 6 VGND
port 2 nsew ground bidirectional
rlabel metal5 s 1056 12672 12836 12992 6 VGND
port 2 nsew ground bidirectional
rlabel metal4 s 2404 2128 2724 13648 6 VPWR
port 3 nsew power bidirectional
rlabel metal4 s 5325 2128 5645 13648 6 VPWR
port 3 nsew power bidirectional
rlabel metal4 s 8246 2128 8566 13648 6 VPWR
port 3 nsew power bidirectional
rlabel metal4 s 11167 2128 11487 13648 6 VPWR
port 3 nsew power bidirectional
rlabel metal5 s 1056 3444 12836 3764 6 VPWR
port 3 nsew power bidirectional
rlabel metal5 s 1056 6300 12836 6620 6 VPWR
port 3 nsew power bidirectional
rlabel metal5 s 1056 9156 12836 9476 6 VPWR
port 3 nsew power bidirectional
rlabel metal5 s 1056 12012 12836 12332 6 VPWR
port 3 nsew power bidirectional
rlabel metal3 s 0 14968 800 15088 6 clk
port 4 nsew signal input
rlabel metal2 s 13542 15266 13598 16066 6 decrease_duty
port 5 nsew signal input
rlabel metal3 s 13122 688 13922 808 6 increase_duty
port 6 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 13922 16066
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 763886
string GDS_FILE /home/veda/Pulse-width-modulator/openlane/pes_pwm/runs/23_11_25_11_08/results/signoff/pes_pwm.magic.gds
string GDS_START 320820
<< end >>

