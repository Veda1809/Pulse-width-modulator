magic
tech sky130A
magscale 1 2
timestamp 1700890849
<< viali >>
rect 5917 13413 5951 13447
rect 4905 13277 4939 13311
rect 5641 13277 5675 13311
rect 5733 13277 5767 13311
rect 5825 13277 5859 13311
rect 6469 13277 6503 13311
rect 6745 13277 6779 13311
rect 12449 13277 12483 13311
rect 12265 13141 12299 13175
rect 6009 12937 6043 12971
rect 4896 12869 4930 12903
rect 6736 12801 6770 12835
rect 7941 12801 7975 12835
rect 8125 12801 8159 12835
rect 4629 12733 4663 12767
rect 6469 12733 6503 12767
rect 7849 12665 7883 12699
rect 4537 12597 4571 12631
rect 8125 12597 8159 12631
rect 5733 12393 5767 12427
rect 7205 12393 7239 12427
rect 4353 12257 4387 12291
rect 8033 12257 8067 12291
rect 4609 12189 4643 12223
rect 5825 12189 5859 12223
rect 7297 12189 7331 12223
rect 7665 12189 7699 12223
rect 8125 12189 8159 12223
rect 8677 12189 8711 12223
rect 6092 12121 6126 12155
rect 6469 11849 6503 11883
rect 8585 11849 8619 11883
rect 8769 11849 8803 11883
rect 4813 11713 4847 11747
rect 5069 11713 5103 11747
rect 6377 11713 6411 11747
rect 6561 11713 6595 11747
rect 7113 11713 7147 11747
rect 7461 11713 7495 11747
rect 8677 11713 8711 11747
rect 8861 11713 8895 11747
rect 4721 11645 4755 11679
rect 7205 11645 7239 11679
rect 6193 11577 6227 11611
rect 6837 11509 6871 11543
rect 6377 11305 6411 11339
rect 8309 11305 8343 11339
rect 4997 11169 5031 11203
rect 5264 11101 5298 11135
rect 6929 11101 6963 11135
rect 7185 11101 7219 11135
rect 3801 10625 3835 10659
rect 4068 10625 4102 10659
rect 3525 10421 3559 10455
rect 5181 10421 5215 10455
rect 5733 10421 5767 10455
rect 4077 10217 4111 10251
rect 2237 10013 2271 10047
rect 4721 10013 4755 10047
rect 4813 10013 4847 10047
rect 5089 10013 5123 10047
rect 5181 10013 5215 10047
rect 6653 10013 6687 10047
rect 2504 9945 2538 9979
rect 4537 9945 4571 9979
rect 5448 9945 5482 9979
rect 6920 9945 6954 9979
rect 3617 9877 3651 9911
rect 4813 9877 4847 9911
rect 6561 9877 6595 9911
rect 8033 9877 8067 9911
rect 4721 9673 4755 9707
rect 5080 9605 5114 9639
rect 3341 9537 3375 9571
rect 3608 9537 3642 9571
rect 4813 9537 4847 9571
rect 6377 9537 6411 9571
rect 6929 9537 6963 9571
rect 7389 9537 7423 9571
rect 7481 9537 7515 9571
rect 2789 9469 2823 9503
rect 7205 9469 7239 9503
rect 6193 9333 6227 9367
rect 7481 9333 7515 9367
rect 6837 9129 6871 9163
rect 3801 8993 3835 9027
rect 1869 8925 1903 8959
rect 2145 8925 2179 8959
rect 3617 8925 3651 8959
rect 4057 8925 4091 8959
rect 5457 8925 5491 8959
rect 6929 8925 6963 8959
rect 7205 8925 7239 8959
rect 7665 8925 7699 8959
rect 7941 8925 7975 8959
rect 8309 8925 8343 8959
rect 8953 8925 8987 8959
rect 9229 8925 9263 8959
rect 5724 8857 5758 8891
rect 7757 8857 7791 8891
rect 5181 8789 5215 8823
rect 3433 8585 3467 8619
rect 4997 8585 5031 8619
rect 7757 8585 7791 8619
rect 7941 8585 7975 8619
rect 9965 8585 9999 8619
rect 1860 8517 1894 8551
rect 5089 8517 5123 8551
rect 5273 8517 5307 8551
rect 5733 8517 5767 8551
rect 6644 8517 6678 8551
rect 8668 8517 8702 8551
rect 3249 8449 3283 8483
rect 3341 8449 3375 8483
rect 3525 8449 3559 8483
rect 3801 8449 3835 8483
rect 3893 8449 3927 8483
rect 3985 8449 4019 8483
rect 4353 8449 4387 8483
rect 4629 8449 4663 8483
rect 4905 8449 4939 8483
rect 6009 8449 6043 8483
rect 6193 8449 6227 8483
rect 7849 8449 7883 8483
rect 8033 8449 8067 8483
rect 9873 8449 9907 8483
rect 10057 8449 10091 8483
rect 1593 8381 1627 8415
rect 3617 8381 3651 8415
rect 6101 8381 6135 8415
rect 6377 8381 6411 8415
rect 8401 8381 8435 8415
rect 2973 8313 3007 8347
rect 3893 8313 3927 8347
rect 4721 8313 4755 8347
rect 5365 8313 5399 8347
rect 9781 8313 9815 8347
rect 4077 8245 4111 8279
rect 5733 8245 5767 8279
rect 5917 8245 5951 8279
rect 2789 8041 2823 8075
rect 10333 8041 10367 8075
rect 1409 7905 1443 7939
rect 5733 7905 5767 7939
rect 8953 7905 8987 7939
rect 1676 7837 1710 7871
rect 3893 7837 3927 7871
rect 4077 7837 4111 7871
rect 4537 7837 4571 7871
rect 5825 7837 5859 7871
rect 7849 7837 7883 7871
rect 8125 7837 8159 7871
rect 3985 7769 4019 7803
rect 7665 7769 7699 7803
rect 9220 7769 9254 7803
rect 4445 7701 4479 7735
rect 5089 7701 5123 7735
rect 7113 7701 7147 7735
rect 5825 7497 5859 7531
rect 7757 7497 7791 7531
rect 10977 7497 11011 7531
rect 2605 7429 2639 7463
rect 4353 7429 4387 7463
rect 6644 7429 6678 7463
rect 9036 7429 9070 7463
rect 4701 7361 4735 7395
rect 6009 7361 6043 7395
rect 6377 7361 6411 7395
rect 7941 7361 7975 7395
rect 8125 7361 8159 7395
rect 8309 7361 8343 7395
rect 8493 7361 8527 7395
rect 10241 7361 10275 7395
rect 11161 7361 11195 7395
rect 4445 7293 4479 7327
rect 8677 7293 8711 7327
rect 8769 7293 8803 7327
rect 10793 7293 10827 7327
rect 2237 7157 2271 7191
rect 2513 7157 2547 7191
rect 6193 7157 6227 7191
rect 10149 7157 10183 7191
rect 3617 6953 3651 6987
rect 3893 6953 3927 6987
rect 6561 6953 6595 6987
rect 7113 6885 7147 6919
rect 3801 6817 3835 6851
rect 3985 6817 4019 6851
rect 8493 6817 8527 6851
rect 9321 6817 9355 6851
rect 9505 6817 9539 6851
rect 1961 6749 1995 6783
rect 2237 6749 2271 6783
rect 4353 6749 4387 6783
rect 4629 6749 4663 6783
rect 4813 6749 4847 6783
rect 4997 6749 5031 6783
rect 5181 6749 5215 6783
rect 5275 6749 5309 6783
rect 8226 6749 8260 6783
rect 8769 6749 8803 6783
rect 9597 6749 9631 6783
rect 2482 6681 2516 6715
rect 4169 6681 4203 6715
rect 4077 6613 4111 6647
rect 8677 6613 8711 6647
rect 9965 6613 9999 6647
rect 1869 6409 1903 6443
rect 3433 6409 3467 6443
rect 7113 6409 7147 6443
rect 9137 6409 9171 6443
rect 10241 6409 10275 6443
rect 2298 6341 2332 6375
rect 4712 6341 4746 6375
rect 6009 6341 6043 6375
rect 10149 6341 10183 6375
rect 1777 6273 1811 6307
rect 1961 6273 1995 6307
rect 3525 6273 3559 6307
rect 3709 6273 3743 6307
rect 3801 6273 3835 6307
rect 3893 6273 3927 6307
rect 4077 6273 4111 6307
rect 4169 6273 4203 6307
rect 4445 6273 4479 6307
rect 5917 6273 5951 6307
rect 6193 6273 6227 6307
rect 7021 6273 7055 6307
rect 7389 6273 7423 6307
rect 7757 6273 7791 6307
rect 8125 6273 8159 6307
rect 8769 6273 8803 6307
rect 9045 6273 9079 6307
rect 9321 6273 9355 6307
rect 10425 6273 10459 6307
rect 10793 6273 10827 6307
rect 11253 6273 11287 6307
rect 2053 6205 2087 6239
rect 4261 6205 4295 6239
rect 6377 6205 6411 6239
rect 7297 6205 7331 6239
rect 8217 6205 8251 6239
rect 8677 6205 8711 6239
rect 9505 6205 9539 6239
rect 10701 6205 10735 6239
rect 10885 6205 10919 6239
rect 5825 6137 5859 6171
rect 6101 6137 6135 6171
rect 8493 6137 8527 6171
rect 1685 6069 1719 6103
rect 3801 6069 3835 6103
rect 4353 6069 4387 6103
rect 10609 6069 10643 6103
rect 11069 6069 11103 6103
rect 3617 5865 3651 5899
rect 5457 5865 5491 5899
rect 8033 5865 8067 5899
rect 6009 5729 6043 5763
rect 7389 5729 7423 5763
rect 8217 5729 8251 5763
rect 8401 5729 8435 5763
rect 9045 5729 9079 5763
rect 11069 5729 11103 5763
rect 1961 5661 1995 5695
rect 2145 5661 2179 5695
rect 2237 5661 2271 5695
rect 3801 5661 3835 5695
rect 5273 5661 5307 5695
rect 5365 5661 5399 5695
rect 5641 5661 5675 5695
rect 5825 5661 5859 5695
rect 6101 5661 6135 5695
rect 6469 5661 6503 5695
rect 6653 5661 6687 5695
rect 7297 5661 7331 5695
rect 7757 5661 7791 5695
rect 7960 5661 7994 5695
rect 8125 5661 8159 5695
rect 8309 5661 8343 5695
rect 9312 5661 9346 5695
rect 11437 5661 11471 5695
rect 2482 5593 2516 5627
rect 4046 5593 4080 5627
rect 5549 5593 5583 5627
rect 8585 5593 8619 5627
rect 1961 5525 1995 5559
rect 5181 5525 5215 5559
rect 6653 5525 6687 5559
rect 7849 5525 7883 5559
rect 8493 5525 8527 5559
rect 10425 5525 10459 5559
rect 10517 5525 10551 5559
rect 11253 5525 11287 5559
rect 6561 5321 6595 5355
rect 6653 5321 6687 5355
rect 9413 5321 9447 5355
rect 9781 5321 9815 5355
rect 4353 5253 4387 5287
rect 10333 5253 10367 5287
rect 1869 5185 1903 5219
rect 2237 5185 2271 5219
rect 2421 5185 2455 5219
rect 2513 5185 2547 5219
rect 5650 5185 5684 5219
rect 6009 5185 6043 5219
rect 6193 5185 6227 5219
rect 6729 5207 6763 5241
rect 7021 5185 7055 5219
rect 7297 5185 7331 5219
rect 7665 5185 7699 5219
rect 7849 5185 7883 5219
rect 8125 5185 8159 5219
rect 8493 5185 8527 5219
rect 8769 5185 8803 5219
rect 8953 5185 8987 5219
rect 10425 5183 10459 5217
rect 2789 5117 2823 5151
rect 5917 5117 5951 5151
rect 6377 5117 6411 5151
rect 6837 5117 6871 5151
rect 9873 5117 9907 5151
rect 9965 5117 9999 5151
rect 7113 5049 7147 5083
rect 7205 5049 7239 5083
rect 8585 5049 8619 5083
rect 1685 4981 1719 5015
rect 2053 4981 2087 5015
rect 4537 4981 4571 5015
rect 6101 4981 6135 5015
rect 6653 4981 6687 5015
rect 7757 4981 7791 5015
rect 4721 4777 4755 4811
rect 9781 4777 9815 4811
rect 9873 4777 9907 4811
rect 3801 4709 3835 4743
rect 4905 4709 4939 4743
rect 2973 4641 3007 4675
rect 4997 4641 5031 4675
rect 5457 4641 5491 4675
rect 6009 4641 6043 4675
rect 8033 4641 8067 4675
rect 9137 4641 9171 4675
rect 9229 4641 9263 4675
rect 9781 4641 9815 4675
rect 1409 4573 1443 4607
rect 3617 4573 3651 4607
rect 4353 4573 4387 4607
rect 5181 4573 5215 4607
rect 5273 4573 5307 4607
rect 5365 4573 5399 4607
rect 5641 4573 5675 4607
rect 5733 4573 5767 4607
rect 6193 4573 6227 4607
rect 6285 4573 6319 4607
rect 6561 4573 6595 4607
rect 6929 4573 6963 4607
rect 7481 4573 7515 4607
rect 7757 4573 7791 4607
rect 8125 4573 8159 4607
rect 8769 4573 8803 4607
rect 9312 4573 9346 4607
rect 9413 4573 9447 4607
rect 9965 4573 9999 4607
rect 10241 4573 10275 4607
rect 1676 4505 1710 4539
rect 4537 4505 4571 4539
rect 6469 4505 6503 4539
rect 9597 4505 9631 4539
rect 2789 4437 2823 4471
rect 4747 4437 4781 4471
rect 5825 4437 5859 4471
rect 6009 4437 6043 4471
rect 8953 4437 8987 4471
rect 10057 4437 10091 4471
rect 3065 4233 3099 4267
rect 3893 4233 3927 4267
rect 5089 4233 5123 4267
rect 5457 4233 5491 4267
rect 8953 4233 8987 4267
rect 9045 4233 9079 4267
rect 2706 4165 2740 4199
rect 3249 4165 3283 4199
rect 3709 4165 3743 4199
rect 5825 4165 5859 4199
rect 2973 4097 3007 4131
rect 3969 4097 4003 4131
rect 4077 4097 4111 4131
rect 4261 4097 4295 4131
rect 4353 4097 4387 4131
rect 4445 4097 4479 4131
rect 4721 4097 4755 4131
rect 4813 4097 4847 4131
rect 4997 4097 5031 4131
rect 5273 4097 5307 4131
rect 5549 4097 5583 4131
rect 5641 4097 5675 4131
rect 5917 4097 5951 4131
rect 6009 4097 6043 4131
rect 6633 4097 6667 4131
rect 8125 4097 8159 4131
rect 8217 4097 8251 4131
rect 8585 4097 8619 4131
rect 8677 4097 8711 4131
rect 8769 4097 8803 4131
rect 9137 4097 9171 4131
rect 9496 4097 9530 4131
rect 3617 4029 3651 4063
rect 6377 4029 6411 4063
rect 9229 4029 9263 4063
rect 3709 3961 3743 3995
rect 8861 3961 8895 3995
rect 1593 3893 1627 3927
rect 3249 3893 3283 3927
rect 4629 3893 4663 3927
rect 4997 3893 5031 3927
rect 6193 3893 6227 3927
rect 7757 3893 7791 3927
rect 8309 3893 8343 3927
rect 10609 3893 10643 3927
rect 7113 3689 7147 3723
rect 9045 3689 9079 3723
rect 9413 3689 9447 3723
rect 10425 3689 10459 3723
rect 1409 3621 1443 3655
rect 2789 3553 2823 3587
rect 4169 3553 4203 3587
rect 7021 3553 7055 3587
rect 9781 3553 9815 3587
rect 3433 3485 3467 3519
rect 3985 3485 4019 3519
rect 4077 3485 4111 3519
rect 4261 3485 4295 3519
rect 4445 3485 4479 3519
rect 4721 3485 4755 3519
rect 4837 3485 4871 3519
rect 5273 3485 5307 3519
rect 7665 3485 7699 3519
rect 8493 3485 8527 3519
rect 8953 3485 8987 3519
rect 9229 3485 9263 3519
rect 9965 3485 9999 3519
rect 2544 3417 2578 3451
rect 2881 3417 2915 3451
rect 4629 3417 4663 3451
rect 10057 3417 10091 3451
rect 3801 3349 3835 3383
rect 4997 3349 5031 3383
rect 7941 3349 7975 3383
rect 1869 3145 1903 3179
rect 6101 3145 6135 3179
rect 6469 3145 6503 3179
rect 7665 3145 7699 3179
rect 9413 3145 9447 3179
rect 1593 3077 1627 3111
rect 1777 3077 1811 3111
rect 1501 3009 1535 3043
rect 2053 3009 2087 3043
rect 2237 3009 2271 3043
rect 3065 3009 3099 3043
rect 4721 3009 4755 3043
rect 5089 3009 5123 3043
rect 5273 3009 5307 3043
rect 5549 3009 5583 3043
rect 6009 3009 6043 3043
rect 6377 3009 6411 3043
rect 6653 3009 6687 3043
rect 7205 3009 7239 3043
rect 7389 3009 7423 3043
rect 7757 3009 7791 3043
rect 7849 3009 7883 3043
rect 2329 2941 2363 2975
rect 3709 2941 3743 2975
rect 3801 2941 3835 2975
rect 4905 2941 4939 2975
rect 4997 2941 5031 2975
rect 5641 2941 5675 2975
rect 5917 2941 5951 2975
rect 6837 2941 6871 2975
rect 7297 2941 7331 2975
rect 8125 2941 8159 2975
rect 1777 2873 1811 2907
rect 6745 2873 6779 2907
rect 7021 2873 7055 2907
rect 2973 2805 3007 2839
rect 4445 2805 4479 2839
rect 4537 2805 4571 2839
rect 6837 2805 6871 2839
rect 2145 2601 2179 2635
rect 2789 2601 2823 2635
rect 6469 2601 6503 2635
rect 8125 2601 8159 2635
rect 8585 2601 8619 2635
rect 8677 2601 8711 2635
rect 9045 2601 9079 2635
rect 12265 2601 12299 2635
rect 2237 2465 2271 2499
rect 2605 2465 2639 2499
rect 5181 2465 5215 2499
rect 6745 2465 6779 2499
rect 8493 2465 8527 2499
rect 2150 2397 2184 2431
rect 3065 2397 3099 2431
rect 3341 2397 3375 2431
rect 3617 2397 3651 2431
rect 4914 2397 4948 2431
rect 5641 2397 5675 2431
rect 5825 2397 5859 2431
rect 6377 2397 6411 2431
rect 7001 2397 7035 2431
rect 8769 2397 8803 2431
rect 8953 2397 8987 2431
rect 9137 2397 9171 2431
rect 12449 2397 12483 2431
rect 1409 2329 1443 2363
rect 1777 2329 1811 2363
rect 3157 2329 3191 2363
rect 3525 2329 3559 2363
rect 5457 2329 5491 2363
rect 2513 2261 2547 2295
rect 2973 2261 3007 2295
rect 3801 2261 3835 2295
rect 5273 2261 5307 2295
rect 5917 2261 5951 2295
<< metal1 >>
rect 4062 13812 4068 13864
rect 4120 13852 4126 13864
rect 5810 13852 5816 13864
rect 4120 13824 5816 13852
rect 4120 13812 4126 13824
rect 5810 13812 5816 13824
rect 5868 13812 5874 13864
rect 1104 13626 12788 13648
rect 1104 13574 2410 13626
rect 2462 13574 2474 13626
rect 2526 13574 2538 13626
rect 2590 13574 2602 13626
rect 2654 13574 2666 13626
rect 2718 13574 5331 13626
rect 5383 13574 5395 13626
rect 5447 13574 5459 13626
rect 5511 13574 5523 13626
rect 5575 13574 5587 13626
rect 5639 13574 8252 13626
rect 8304 13574 8316 13626
rect 8368 13574 8380 13626
rect 8432 13574 8444 13626
rect 8496 13574 8508 13626
rect 8560 13574 11173 13626
rect 11225 13574 11237 13626
rect 11289 13574 11301 13626
rect 11353 13574 11365 13626
rect 11417 13574 11429 13626
rect 11481 13574 12788 13626
rect 1104 13552 12788 13574
rect 5905 13447 5963 13453
rect 5905 13413 5917 13447
rect 5951 13444 5963 13447
rect 6546 13444 6552 13456
rect 5951 13416 6552 13444
rect 5951 13413 5963 13416
rect 5905 13407 5963 13413
rect 6546 13404 6552 13416
rect 6604 13404 6610 13456
rect 7282 13376 7288 13388
rect 5736 13348 7288 13376
rect 4890 13268 4896 13320
rect 4948 13268 4954 13320
rect 5626 13268 5632 13320
rect 5684 13268 5690 13320
rect 5736 13317 5764 13348
rect 7282 13336 7288 13348
rect 7340 13336 7346 13388
rect 13538 13376 13544 13388
rect 12452 13348 13544 13376
rect 5721 13311 5779 13317
rect 5721 13277 5733 13311
rect 5767 13277 5779 13311
rect 5721 13271 5779 13277
rect 5813 13311 5871 13317
rect 5813 13277 5825 13311
rect 5859 13277 5871 13311
rect 5813 13271 5871 13277
rect 5828 13172 5856 13271
rect 6454 13268 6460 13320
rect 6512 13268 6518 13320
rect 6730 13268 6736 13320
rect 6788 13268 6794 13320
rect 12452 13317 12480 13348
rect 13538 13336 13544 13348
rect 13596 13336 13602 13388
rect 12437 13311 12495 13317
rect 12437 13277 12449 13311
rect 12483 13277 12495 13311
rect 12437 13271 12495 13277
rect 5902 13172 5908 13184
rect 5828 13144 5908 13172
rect 5902 13132 5908 13144
rect 5960 13132 5966 13184
rect 12250 13132 12256 13184
rect 12308 13132 12314 13184
rect 1104 13082 12788 13104
rect 1104 13030 3070 13082
rect 3122 13030 3134 13082
rect 3186 13030 3198 13082
rect 3250 13030 3262 13082
rect 3314 13030 3326 13082
rect 3378 13030 5991 13082
rect 6043 13030 6055 13082
rect 6107 13030 6119 13082
rect 6171 13030 6183 13082
rect 6235 13030 6247 13082
rect 6299 13030 8912 13082
rect 8964 13030 8976 13082
rect 9028 13030 9040 13082
rect 9092 13030 9104 13082
rect 9156 13030 9168 13082
rect 9220 13030 11833 13082
rect 11885 13030 11897 13082
rect 11949 13030 11961 13082
rect 12013 13030 12025 13082
rect 12077 13030 12089 13082
rect 12141 13030 12788 13082
rect 1104 13008 12788 13030
rect 5902 12928 5908 12980
rect 5960 12968 5966 12980
rect 5997 12971 6055 12977
rect 5997 12968 6009 12971
rect 5960 12940 6009 12968
rect 5960 12928 5966 12940
rect 5997 12937 6009 12940
rect 6043 12937 6055 12971
rect 5997 12931 6055 12937
rect 4890 12909 4896 12912
rect 4884 12900 4896 12909
rect 4851 12872 4896 12900
rect 4884 12863 4896 12872
rect 4890 12860 4896 12863
rect 4948 12860 4954 12912
rect 6730 12841 6736 12844
rect 6724 12832 6736 12841
rect 6691 12804 6736 12832
rect 6724 12795 6736 12804
rect 6730 12792 6736 12795
rect 6788 12792 6794 12844
rect 7926 12792 7932 12844
rect 7984 12792 7990 12844
rect 8113 12835 8171 12841
rect 8113 12801 8125 12835
rect 8159 12801 8171 12835
rect 8113 12795 8171 12801
rect 4614 12724 4620 12776
rect 4672 12724 4678 12776
rect 6454 12724 6460 12776
rect 6512 12724 6518 12776
rect 8128 12764 8156 12795
rect 7852 12736 8156 12764
rect 7852 12705 7880 12736
rect 7837 12699 7895 12705
rect 7837 12665 7849 12699
rect 7883 12665 7895 12699
rect 7837 12659 7895 12665
rect 4522 12588 4528 12640
rect 4580 12588 4586 12640
rect 8110 12588 8116 12640
rect 8168 12588 8174 12640
rect 1104 12538 12788 12560
rect 1104 12486 2410 12538
rect 2462 12486 2474 12538
rect 2526 12486 2538 12538
rect 2590 12486 2602 12538
rect 2654 12486 2666 12538
rect 2718 12486 5331 12538
rect 5383 12486 5395 12538
rect 5447 12486 5459 12538
rect 5511 12486 5523 12538
rect 5575 12486 5587 12538
rect 5639 12486 8252 12538
rect 8304 12486 8316 12538
rect 8368 12486 8380 12538
rect 8432 12486 8444 12538
rect 8496 12486 8508 12538
rect 8560 12486 11173 12538
rect 11225 12486 11237 12538
rect 11289 12486 11301 12538
rect 11353 12486 11365 12538
rect 11417 12486 11429 12538
rect 11481 12486 12788 12538
rect 1104 12464 12788 12486
rect 4614 12424 4620 12436
rect 4356 12396 4620 12424
rect 4356 12297 4384 12396
rect 4614 12384 4620 12396
rect 4672 12384 4678 12436
rect 5718 12384 5724 12436
rect 5776 12384 5782 12436
rect 7193 12427 7251 12433
rect 7193 12393 7205 12427
rect 7239 12424 7251 12427
rect 7926 12424 7932 12436
rect 7239 12396 7932 12424
rect 7239 12393 7251 12396
rect 7193 12387 7251 12393
rect 7926 12384 7932 12396
rect 7984 12384 7990 12436
rect 4341 12291 4399 12297
rect 4341 12257 4353 12291
rect 4387 12257 4399 12291
rect 4341 12251 4399 12257
rect 8018 12248 8024 12300
rect 8076 12248 8082 12300
rect 4430 12180 4436 12232
rect 4488 12220 4494 12232
rect 4597 12223 4655 12229
rect 4597 12220 4609 12223
rect 4488 12192 4609 12220
rect 4488 12180 4494 12192
rect 4597 12189 4609 12192
rect 4643 12189 4655 12223
rect 4597 12183 4655 12189
rect 5813 12223 5871 12229
rect 5813 12189 5825 12223
rect 5859 12220 5871 12223
rect 6454 12220 6460 12232
rect 5859 12192 6460 12220
rect 5859 12189 5871 12192
rect 5813 12183 5871 12189
rect 6454 12180 6460 12192
rect 6512 12220 6518 12232
rect 6822 12220 6828 12232
rect 6512 12192 6828 12220
rect 6512 12180 6518 12192
rect 6822 12180 6828 12192
rect 6880 12180 6886 12232
rect 7282 12180 7288 12232
rect 7340 12180 7346 12232
rect 7650 12180 7656 12232
rect 7708 12180 7714 12232
rect 8110 12180 8116 12232
rect 8168 12180 8174 12232
rect 8662 12180 8668 12232
rect 8720 12180 8726 12232
rect 6080 12155 6138 12161
rect 6080 12121 6092 12155
rect 6126 12152 6138 12155
rect 6362 12152 6368 12164
rect 6126 12124 6368 12152
rect 6126 12121 6138 12124
rect 6080 12115 6138 12121
rect 6362 12112 6368 12124
rect 6420 12112 6426 12164
rect 1104 11994 12788 12016
rect 1104 11942 3070 11994
rect 3122 11942 3134 11994
rect 3186 11942 3198 11994
rect 3250 11942 3262 11994
rect 3314 11942 3326 11994
rect 3378 11942 5991 11994
rect 6043 11942 6055 11994
rect 6107 11942 6119 11994
rect 6171 11942 6183 11994
rect 6235 11942 6247 11994
rect 6299 11942 8912 11994
rect 8964 11942 8976 11994
rect 9028 11942 9040 11994
rect 9092 11942 9104 11994
rect 9156 11942 9168 11994
rect 9220 11942 11833 11994
rect 11885 11942 11897 11994
rect 11949 11942 11961 11994
rect 12013 11942 12025 11994
rect 12077 11942 12089 11994
rect 12141 11942 12788 11994
rect 1104 11920 12788 11942
rect 6457 11883 6515 11889
rect 6457 11849 6469 11883
rect 6503 11880 6515 11883
rect 7650 11880 7656 11892
rect 6503 11852 7656 11880
rect 6503 11849 6515 11852
rect 6457 11843 6515 11849
rect 7650 11840 7656 11852
rect 7708 11840 7714 11892
rect 8573 11883 8631 11889
rect 8573 11849 8585 11883
rect 8619 11849 8631 11883
rect 8573 11843 8631 11849
rect 4614 11704 4620 11756
rect 4672 11744 4678 11756
rect 4801 11747 4859 11753
rect 4801 11744 4813 11747
rect 4672 11716 4813 11744
rect 4672 11704 4678 11716
rect 4801 11713 4813 11716
rect 4847 11713 4859 11747
rect 5057 11747 5115 11753
rect 5057 11744 5069 11747
rect 4801 11707 4859 11713
rect 4899 11716 5069 11744
rect 4709 11679 4767 11685
rect 4709 11645 4721 11679
rect 4755 11676 4767 11679
rect 4899 11676 4927 11716
rect 5057 11713 5069 11716
rect 5103 11713 5115 11747
rect 5057 11707 5115 11713
rect 6362 11704 6368 11756
rect 6420 11704 6426 11756
rect 6549 11747 6607 11753
rect 6549 11713 6561 11747
rect 6595 11713 6607 11747
rect 6549 11707 6607 11713
rect 7101 11747 7159 11753
rect 7101 11713 7113 11747
rect 7147 11744 7159 11747
rect 7449 11747 7507 11753
rect 7449 11744 7461 11747
rect 7147 11716 7461 11744
rect 7147 11713 7159 11716
rect 7101 11707 7159 11713
rect 7449 11713 7461 11716
rect 7495 11713 7507 11747
rect 8588 11744 8616 11843
rect 8662 11840 8668 11892
rect 8720 11880 8726 11892
rect 8757 11883 8815 11889
rect 8757 11880 8769 11883
rect 8720 11852 8769 11880
rect 8720 11840 8726 11852
rect 8757 11849 8769 11852
rect 8803 11849 8815 11883
rect 8757 11843 8815 11849
rect 8665 11747 8723 11753
rect 8665 11744 8677 11747
rect 8588 11716 8677 11744
rect 7449 11707 7507 11713
rect 8665 11713 8677 11716
rect 8711 11713 8723 11747
rect 8665 11707 8723 11713
rect 6564 11676 6592 11707
rect 8846 11704 8852 11756
rect 8904 11704 8910 11756
rect 4755 11648 4927 11676
rect 6196 11648 6592 11676
rect 4755 11645 4767 11648
rect 4709 11639 4767 11645
rect 6196 11617 6224 11648
rect 6822 11636 6828 11688
rect 6880 11676 6886 11688
rect 7193 11679 7251 11685
rect 7193 11676 7205 11679
rect 6880 11648 7205 11676
rect 6880 11636 6886 11648
rect 7193 11645 7205 11648
rect 7239 11645 7251 11679
rect 7193 11639 7251 11645
rect 6181 11611 6239 11617
rect 6181 11577 6193 11611
rect 6227 11577 6239 11611
rect 6181 11571 6239 11577
rect 6825 11543 6883 11549
rect 6825 11509 6837 11543
rect 6871 11540 6883 11543
rect 6914 11540 6920 11552
rect 6871 11512 6920 11540
rect 6871 11509 6883 11512
rect 6825 11503 6883 11509
rect 6914 11500 6920 11512
rect 6972 11500 6978 11552
rect 1104 11450 12788 11472
rect 1104 11398 2410 11450
rect 2462 11398 2474 11450
rect 2526 11398 2538 11450
rect 2590 11398 2602 11450
rect 2654 11398 2666 11450
rect 2718 11398 5331 11450
rect 5383 11398 5395 11450
rect 5447 11398 5459 11450
rect 5511 11398 5523 11450
rect 5575 11398 5587 11450
rect 5639 11398 8252 11450
rect 8304 11398 8316 11450
rect 8368 11398 8380 11450
rect 8432 11398 8444 11450
rect 8496 11398 8508 11450
rect 8560 11398 11173 11450
rect 11225 11398 11237 11450
rect 11289 11398 11301 11450
rect 11353 11398 11365 11450
rect 11417 11398 11429 11450
rect 11481 11398 12788 11450
rect 1104 11376 12788 11398
rect 6362 11296 6368 11348
rect 6420 11296 6426 11348
rect 6914 11296 6920 11348
rect 6972 11296 6978 11348
rect 8297 11339 8355 11345
rect 8297 11305 8309 11339
rect 8343 11336 8355 11339
rect 8846 11336 8852 11348
rect 8343 11308 8852 11336
rect 8343 11305 8355 11308
rect 8297 11299 8355 11305
rect 8846 11296 8852 11308
rect 8904 11296 8910 11348
rect 4614 11160 4620 11212
rect 4672 11200 4678 11212
rect 4985 11203 5043 11209
rect 4985 11200 4997 11203
rect 4672 11172 4997 11200
rect 4672 11160 4678 11172
rect 4985 11169 4997 11172
rect 5031 11169 5043 11203
rect 6546 11200 6552 11212
rect 4985 11163 5043 11169
rect 6288 11172 6552 11200
rect 5252 11135 5310 11141
rect 5252 11101 5264 11135
rect 5298 11132 5310 11135
rect 6288 11132 6316 11172
rect 6546 11160 6552 11172
rect 6604 11160 6610 11212
rect 6932 11200 6960 11296
rect 6932 11172 7052 11200
rect 5298 11104 6316 11132
rect 5298 11101 5310 11104
rect 5252 11095 5310 11101
rect 6362 11092 6368 11144
rect 6420 11132 6426 11144
rect 6822 11132 6828 11144
rect 6420 11104 6828 11132
rect 6420 11092 6426 11104
rect 6822 11092 6828 11104
rect 6880 11132 6886 11144
rect 6917 11135 6975 11141
rect 6917 11132 6929 11135
rect 6880 11104 6929 11132
rect 6880 11092 6886 11104
rect 6917 11101 6929 11104
rect 6963 11101 6975 11135
rect 7024 11132 7052 11172
rect 7173 11135 7231 11141
rect 7173 11132 7185 11135
rect 7024 11104 7185 11132
rect 6917 11095 6975 11101
rect 7173 11101 7185 11104
rect 7219 11101 7231 11135
rect 7173 11095 7231 11101
rect 1104 10906 12788 10928
rect 1104 10854 3070 10906
rect 3122 10854 3134 10906
rect 3186 10854 3198 10906
rect 3250 10854 3262 10906
rect 3314 10854 3326 10906
rect 3378 10854 5991 10906
rect 6043 10854 6055 10906
rect 6107 10854 6119 10906
rect 6171 10854 6183 10906
rect 6235 10854 6247 10906
rect 6299 10854 8912 10906
rect 8964 10854 8976 10906
rect 9028 10854 9040 10906
rect 9092 10854 9104 10906
rect 9156 10854 9168 10906
rect 9220 10854 11833 10906
rect 11885 10854 11897 10906
rect 11949 10854 11961 10906
rect 12013 10854 12025 10906
rect 12077 10854 12089 10906
rect 12141 10854 12788 10906
rect 1104 10832 12788 10854
rect 4614 10792 4620 10804
rect 3804 10764 4620 10792
rect 3804 10665 3832 10764
rect 4614 10752 4620 10764
rect 4672 10752 4678 10804
rect 4062 10665 4068 10668
rect 3789 10659 3847 10665
rect 3789 10625 3801 10659
rect 3835 10625 3847 10659
rect 3789 10619 3847 10625
rect 4056 10619 4068 10665
rect 4062 10616 4068 10619
rect 4120 10616 4126 10668
rect 3513 10455 3571 10461
rect 3513 10421 3525 10455
rect 3559 10452 3571 10455
rect 3602 10452 3608 10464
rect 3559 10424 3608 10452
rect 3559 10421 3571 10424
rect 3513 10415 3571 10421
rect 3602 10412 3608 10424
rect 3660 10412 3666 10464
rect 5166 10412 5172 10464
rect 5224 10412 5230 10464
rect 5718 10412 5724 10464
rect 5776 10412 5782 10464
rect 1104 10362 12788 10384
rect 1104 10310 2410 10362
rect 2462 10310 2474 10362
rect 2526 10310 2538 10362
rect 2590 10310 2602 10362
rect 2654 10310 2666 10362
rect 2718 10310 5331 10362
rect 5383 10310 5395 10362
rect 5447 10310 5459 10362
rect 5511 10310 5523 10362
rect 5575 10310 5587 10362
rect 5639 10310 8252 10362
rect 8304 10310 8316 10362
rect 8368 10310 8380 10362
rect 8432 10310 8444 10362
rect 8496 10310 8508 10362
rect 8560 10310 11173 10362
rect 11225 10310 11237 10362
rect 11289 10310 11301 10362
rect 11353 10310 11365 10362
rect 11417 10310 11429 10362
rect 11481 10310 12788 10362
rect 1104 10288 12788 10310
rect 4062 10208 4068 10260
rect 4120 10208 4126 10260
rect 5166 10208 5172 10260
rect 5224 10208 5230 10260
rect 5184 10112 5212 10208
rect 4816 10084 5212 10112
rect 1394 10004 1400 10056
rect 1452 10044 1458 10056
rect 2225 10047 2283 10053
rect 2225 10044 2237 10047
rect 1452 10016 2237 10044
rect 1452 10004 1458 10016
rect 2225 10013 2237 10016
rect 2271 10013 2283 10047
rect 2225 10007 2283 10013
rect 4706 10004 4712 10056
rect 4764 10004 4770 10056
rect 4816 10053 4844 10084
rect 4801 10047 4859 10053
rect 4801 10013 4813 10047
rect 4847 10013 4859 10047
rect 4801 10007 4859 10013
rect 5074 10004 5080 10056
rect 5132 10004 5138 10056
rect 5169 10047 5227 10053
rect 5169 10013 5181 10047
rect 5215 10044 5227 10047
rect 6362 10044 6368 10056
rect 5215 10016 6368 10044
rect 5215 10013 5227 10016
rect 5169 10007 5227 10013
rect 6362 10004 6368 10016
rect 6420 10044 6426 10056
rect 6641 10047 6699 10053
rect 6641 10044 6653 10047
rect 6420 10016 6653 10044
rect 6420 10004 6426 10016
rect 6641 10013 6653 10016
rect 6687 10013 6699 10047
rect 6641 10007 6699 10013
rect 2492 9979 2550 9985
rect 2492 9945 2504 9979
rect 2538 9976 2550 9979
rect 2774 9976 2780 9988
rect 2538 9948 2780 9976
rect 2538 9945 2550 9948
rect 2492 9939 2550 9945
rect 2774 9936 2780 9948
rect 2832 9936 2838 9988
rect 4525 9979 4583 9985
rect 4525 9976 4537 9979
rect 3620 9948 4537 9976
rect 3620 9917 3648 9948
rect 4525 9945 4537 9948
rect 4571 9945 4583 9979
rect 4525 9939 4583 9945
rect 5436 9979 5494 9985
rect 5436 9945 5448 9979
rect 5482 9976 5494 9979
rect 5902 9976 5908 9988
rect 5482 9948 5908 9976
rect 5482 9945 5494 9948
rect 5436 9939 5494 9945
rect 5902 9936 5908 9948
rect 5960 9936 5966 9988
rect 6914 9985 6920 9988
rect 6908 9939 6920 9985
rect 6914 9936 6920 9939
rect 6972 9936 6978 9988
rect 3605 9911 3663 9917
rect 3605 9877 3617 9911
rect 3651 9877 3663 9911
rect 3605 9871 3663 9877
rect 4798 9868 4804 9920
rect 4856 9868 4862 9920
rect 6549 9911 6607 9917
rect 6549 9877 6561 9911
rect 6595 9908 6607 9911
rect 7374 9908 7380 9920
rect 6595 9880 7380 9908
rect 6595 9877 6607 9880
rect 6549 9871 6607 9877
rect 7374 9868 7380 9880
rect 7432 9868 7438 9920
rect 8018 9868 8024 9920
rect 8076 9868 8082 9920
rect 1104 9818 12788 9840
rect 1104 9766 3070 9818
rect 3122 9766 3134 9818
rect 3186 9766 3198 9818
rect 3250 9766 3262 9818
rect 3314 9766 3326 9818
rect 3378 9766 5991 9818
rect 6043 9766 6055 9818
rect 6107 9766 6119 9818
rect 6171 9766 6183 9818
rect 6235 9766 6247 9818
rect 6299 9766 8912 9818
rect 8964 9766 8976 9818
rect 9028 9766 9040 9818
rect 9092 9766 9104 9818
rect 9156 9766 9168 9818
rect 9220 9766 11833 9818
rect 11885 9766 11897 9818
rect 11949 9766 11961 9818
rect 12013 9766 12025 9818
rect 12077 9766 12089 9818
rect 12141 9766 12788 9818
rect 1104 9744 12788 9766
rect 4706 9664 4712 9716
rect 4764 9664 4770 9716
rect 8018 9664 8024 9716
rect 8076 9664 8082 9716
rect 3786 9636 3792 9648
rect 3344 9608 3792 9636
rect 1394 9528 1400 9580
rect 1452 9568 1458 9580
rect 3344 9577 3372 9608
rect 3786 9596 3792 9608
rect 3844 9636 3850 9648
rect 5074 9645 5080 9648
rect 5068 9636 5080 9645
rect 3844 9608 4660 9636
rect 5035 9608 5080 9636
rect 3844 9596 3850 9608
rect 4632 9580 4660 9608
rect 5068 9599 5080 9608
rect 5074 9596 5080 9599
rect 5132 9596 5138 9648
rect 3602 9577 3608 9580
rect 3329 9571 3387 9577
rect 3329 9568 3341 9571
rect 1452 9540 3341 9568
rect 1452 9528 1458 9540
rect 3329 9537 3341 9540
rect 3375 9537 3387 9571
rect 3596 9568 3608 9577
rect 3563 9540 3608 9568
rect 3329 9531 3387 9537
rect 3596 9531 3608 9540
rect 3602 9528 3608 9531
rect 3660 9528 3666 9580
rect 4614 9528 4620 9580
rect 4672 9568 4678 9580
rect 4801 9571 4859 9577
rect 4801 9568 4813 9571
rect 4672 9540 4813 9568
rect 4672 9528 4678 9540
rect 4801 9537 4813 9540
rect 4847 9537 4859 9571
rect 4801 9531 4859 9537
rect 5902 9528 5908 9580
rect 5960 9568 5966 9580
rect 6365 9571 6423 9577
rect 6365 9568 6377 9571
rect 5960 9540 6377 9568
rect 5960 9528 5966 9540
rect 6365 9537 6377 9540
rect 6411 9537 6423 9571
rect 6365 9531 6423 9537
rect 6914 9528 6920 9580
rect 6972 9528 6978 9580
rect 7374 9528 7380 9580
rect 7432 9528 7438 9580
rect 7469 9571 7527 9577
rect 7469 9537 7481 9571
rect 7515 9568 7527 9571
rect 8036 9568 8064 9664
rect 7515 9540 8064 9568
rect 7515 9537 7527 9540
rect 7469 9531 7527 9537
rect 2774 9460 2780 9512
rect 2832 9460 2838 9512
rect 7190 9460 7196 9512
rect 7248 9460 7254 9512
rect 5902 9324 5908 9376
rect 5960 9364 5966 9376
rect 6181 9367 6239 9373
rect 6181 9364 6193 9367
rect 5960 9336 6193 9364
rect 5960 9324 5966 9336
rect 6181 9333 6193 9336
rect 6227 9333 6239 9367
rect 6181 9327 6239 9333
rect 7466 9324 7472 9376
rect 7524 9324 7530 9376
rect 1104 9274 12788 9296
rect 1104 9222 2410 9274
rect 2462 9222 2474 9274
rect 2526 9222 2538 9274
rect 2590 9222 2602 9274
rect 2654 9222 2666 9274
rect 2718 9222 5331 9274
rect 5383 9222 5395 9274
rect 5447 9222 5459 9274
rect 5511 9222 5523 9274
rect 5575 9222 5587 9274
rect 5639 9222 8252 9274
rect 8304 9222 8316 9274
rect 8368 9222 8380 9274
rect 8432 9222 8444 9274
rect 8496 9222 8508 9274
rect 8560 9222 11173 9274
rect 11225 9222 11237 9274
rect 11289 9222 11301 9274
rect 11353 9222 11365 9274
rect 11417 9222 11429 9274
rect 11481 9222 12788 9274
rect 1104 9200 12788 9222
rect 6825 9163 6883 9169
rect 6825 9129 6837 9163
rect 6871 9160 6883 9163
rect 7190 9160 7196 9172
rect 6871 9132 7196 9160
rect 6871 9129 6883 9132
rect 6825 9123 6883 9129
rect 7190 9120 7196 9132
rect 7248 9120 7254 9172
rect 7466 9120 7472 9172
rect 7524 9120 7530 9172
rect 3786 8984 3792 9036
rect 3844 8984 3850 9036
rect 1854 8916 1860 8968
rect 1912 8916 1918 8968
rect 2130 8916 2136 8968
rect 2188 8916 2194 8968
rect 3605 8959 3663 8965
rect 3605 8925 3617 8959
rect 3651 8956 3663 8959
rect 4045 8959 4103 8965
rect 4045 8956 4057 8959
rect 3651 8928 4057 8956
rect 3651 8925 3663 8928
rect 3605 8919 3663 8925
rect 4045 8925 4057 8928
rect 4091 8925 4103 8959
rect 4045 8919 4103 8925
rect 5445 8959 5503 8965
rect 5445 8925 5457 8959
rect 5491 8956 5503 8959
rect 5491 8928 6408 8956
rect 5491 8925 5503 8928
rect 5445 8919 5503 8925
rect 6380 8900 6408 8928
rect 6914 8916 6920 8968
rect 6972 8916 6978 8968
rect 7190 8916 7196 8968
rect 7248 8916 7254 8968
rect 7484 8956 7512 9120
rect 7653 8959 7711 8965
rect 7653 8956 7665 8959
rect 7484 8928 7665 8956
rect 7653 8925 7665 8928
rect 7699 8925 7711 8959
rect 7653 8919 7711 8925
rect 7926 8916 7932 8968
rect 7984 8916 7990 8968
rect 8297 8959 8355 8965
rect 8297 8925 8309 8959
rect 8343 8925 8355 8959
rect 8297 8919 8355 8925
rect 3878 8848 3884 8900
rect 3936 8888 3942 8900
rect 5350 8888 5356 8900
rect 3936 8860 5356 8888
rect 3936 8848 3942 8860
rect 5350 8848 5356 8860
rect 5408 8848 5414 8900
rect 5718 8897 5724 8900
rect 5712 8888 5724 8897
rect 5679 8860 5724 8888
rect 5712 8851 5724 8860
rect 5718 8848 5724 8851
rect 5776 8848 5782 8900
rect 6362 8848 6368 8900
rect 6420 8848 6426 8900
rect 7742 8848 7748 8900
rect 7800 8848 7806 8900
rect 8312 8888 8340 8919
rect 8754 8916 8760 8968
rect 8812 8956 8818 8968
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 8812 8928 8953 8956
rect 8812 8916 8818 8928
rect 8941 8925 8953 8928
rect 8987 8925 8999 8959
rect 8941 8919 8999 8925
rect 9217 8959 9275 8965
rect 9217 8925 9229 8959
rect 9263 8956 9275 8959
rect 9306 8956 9312 8968
rect 9263 8928 9312 8956
rect 9263 8925 9275 8928
rect 9217 8919 9275 8925
rect 9306 8916 9312 8928
rect 9364 8916 9370 8968
rect 9950 8888 9956 8900
rect 8312 8860 9956 8888
rect 9950 8848 9956 8860
rect 10008 8848 10014 8900
rect 3786 8780 3792 8832
rect 3844 8820 3850 8832
rect 5166 8820 5172 8832
rect 3844 8792 5172 8820
rect 3844 8780 3850 8792
rect 5166 8780 5172 8792
rect 5224 8780 5230 8832
rect 1104 8730 12788 8752
rect 1104 8678 3070 8730
rect 3122 8678 3134 8730
rect 3186 8678 3198 8730
rect 3250 8678 3262 8730
rect 3314 8678 3326 8730
rect 3378 8678 5991 8730
rect 6043 8678 6055 8730
rect 6107 8678 6119 8730
rect 6171 8678 6183 8730
rect 6235 8678 6247 8730
rect 6299 8678 8912 8730
rect 8964 8678 8976 8730
rect 9028 8678 9040 8730
rect 9092 8678 9104 8730
rect 9156 8678 9168 8730
rect 9220 8678 11833 8730
rect 11885 8678 11897 8730
rect 11949 8678 11961 8730
rect 12013 8678 12025 8730
rect 12077 8678 12089 8730
rect 12141 8678 12788 8730
rect 1104 8656 12788 8678
rect 3421 8619 3479 8625
rect 3421 8585 3433 8619
rect 3467 8616 3479 8619
rect 3970 8616 3976 8628
rect 3467 8588 3976 8616
rect 3467 8585 3479 8588
rect 3421 8579 3479 8585
rect 3970 8576 3976 8588
rect 4028 8576 4034 8628
rect 4798 8616 4804 8628
rect 4356 8588 4804 8616
rect 1854 8557 1860 8560
rect 1848 8548 1860 8557
rect 1815 8520 1860 8548
rect 1848 8511 1860 8520
rect 1854 8508 1860 8511
rect 1912 8508 1918 8560
rect 4154 8548 4160 8560
rect 3252 8520 4160 8548
rect 3252 8489 3280 8520
rect 4154 8508 4160 8520
rect 4212 8508 4218 8560
rect 3237 8483 3295 8489
rect 3237 8449 3249 8483
rect 3283 8449 3295 8483
rect 3237 8443 3295 8449
rect 3326 8440 3332 8492
rect 3384 8440 3390 8492
rect 3513 8483 3571 8489
rect 3513 8449 3525 8483
rect 3559 8449 3571 8483
rect 3513 8443 3571 8449
rect 1394 8372 1400 8424
rect 1452 8412 1458 8424
rect 1581 8415 1639 8421
rect 1581 8412 1593 8415
rect 1452 8384 1593 8412
rect 1452 8372 1458 8384
rect 1581 8381 1593 8384
rect 1627 8381 1639 8415
rect 3528 8412 3556 8443
rect 3786 8440 3792 8492
rect 3844 8440 3850 8492
rect 3878 8440 3884 8492
rect 3936 8440 3942 8492
rect 3970 8440 3976 8492
rect 4028 8440 4034 8492
rect 4356 8489 4384 8588
rect 4798 8576 4804 8588
rect 4856 8616 4862 8628
rect 4985 8619 5043 8625
rect 4985 8616 4997 8619
rect 4856 8588 4997 8616
rect 4856 8576 4862 8588
rect 4985 8585 4997 8588
rect 5031 8585 5043 8619
rect 4985 8579 5043 8585
rect 5166 8576 5172 8628
rect 5224 8576 5230 8628
rect 5350 8576 5356 8628
rect 5408 8616 5414 8628
rect 5902 8616 5908 8628
rect 5408 8588 5908 8616
rect 5408 8576 5414 8588
rect 5902 8576 5908 8588
rect 5960 8616 5966 8628
rect 5960 8588 6224 8616
rect 5960 8576 5966 8588
rect 5077 8551 5135 8557
rect 5077 8548 5089 8551
rect 4448 8520 5089 8548
rect 4341 8483 4399 8489
rect 4341 8449 4353 8483
rect 4387 8449 4399 8483
rect 4341 8443 4399 8449
rect 1581 8375 1639 8381
rect 2976 8384 3556 8412
rect 3605 8415 3663 8421
rect 2976 8353 3004 8384
rect 3605 8381 3617 8415
rect 3651 8412 3663 8415
rect 4448 8412 4476 8520
rect 5077 8517 5089 8520
rect 5123 8517 5135 8551
rect 5077 8511 5135 8517
rect 4617 8483 4675 8489
rect 4617 8449 4629 8483
rect 4663 8449 4675 8483
rect 4617 8443 4675 8449
rect 3651 8384 3832 8412
rect 3651 8381 3663 8384
rect 3605 8375 3663 8381
rect 2961 8347 3019 8353
rect 2961 8313 2973 8347
rect 3007 8313 3019 8347
rect 2961 8307 3019 8313
rect 3804 8276 3832 8384
rect 3896 8384 4476 8412
rect 3896 8353 3924 8384
rect 3881 8347 3939 8353
rect 3881 8313 3893 8347
rect 3927 8313 3939 8347
rect 3881 8307 3939 8313
rect 3988 8316 4200 8344
rect 3988 8276 4016 8316
rect 3804 8248 4016 8276
rect 4062 8236 4068 8288
rect 4120 8236 4126 8288
rect 4172 8276 4200 8316
rect 4522 8276 4528 8288
rect 4172 8248 4528 8276
rect 4522 8236 4528 8248
rect 4580 8236 4586 8288
rect 4632 8276 4660 8443
rect 4890 8440 4896 8492
rect 4948 8440 4954 8492
rect 5184 8480 5212 8576
rect 5261 8551 5319 8557
rect 5261 8517 5273 8551
rect 5307 8548 5319 8551
rect 5718 8548 5724 8560
rect 5307 8520 5724 8548
rect 5307 8517 5319 8520
rect 5261 8511 5319 8517
rect 5718 8508 5724 8520
rect 5776 8508 5782 8560
rect 6196 8489 6224 8588
rect 6914 8576 6920 8628
rect 6972 8576 6978 8628
rect 7745 8619 7803 8625
rect 7745 8585 7757 8619
rect 7791 8585 7803 8619
rect 7745 8579 7803 8585
rect 6632 8551 6690 8557
rect 6632 8517 6644 8551
rect 6678 8548 6690 8551
rect 6932 8548 6960 8576
rect 6678 8520 6960 8548
rect 7760 8548 7788 8579
rect 7926 8576 7932 8628
rect 7984 8576 7990 8628
rect 8754 8576 8760 8628
rect 8812 8576 8818 8628
rect 9950 8576 9956 8628
rect 10008 8576 10014 8628
rect 8656 8551 8714 8557
rect 7760 8520 8064 8548
rect 6678 8517 6690 8520
rect 6632 8511 6690 8517
rect 5997 8483 6055 8489
rect 5997 8480 6009 8483
rect 5184 8452 6009 8480
rect 5997 8449 6009 8452
rect 6043 8449 6055 8483
rect 5997 8443 6055 8449
rect 6181 8483 6239 8489
rect 6181 8449 6193 8483
rect 6227 8449 6239 8483
rect 6181 8443 6239 8449
rect 7834 8440 7840 8492
rect 7892 8440 7898 8492
rect 8036 8489 8064 8520
rect 8656 8517 8668 8551
rect 8702 8548 8714 8551
rect 8772 8548 8800 8576
rect 8702 8520 8800 8548
rect 8702 8517 8714 8520
rect 8656 8511 8714 8517
rect 8021 8483 8079 8489
rect 8021 8449 8033 8483
rect 8067 8449 8079 8483
rect 9861 8483 9919 8489
rect 9861 8480 9873 8483
rect 8021 8443 8079 8449
rect 9784 8452 9873 8480
rect 6089 8415 6147 8421
rect 6089 8412 6101 8415
rect 4899 8384 6101 8412
rect 4706 8304 4712 8356
rect 4764 8304 4770 8356
rect 4899 8276 4927 8384
rect 6089 8381 6101 8384
rect 6135 8381 6147 8415
rect 6089 8375 6147 8381
rect 6365 8415 6423 8421
rect 6365 8381 6377 8415
rect 6411 8381 6423 8415
rect 6365 8375 6423 8381
rect 8389 8415 8447 8421
rect 8389 8381 8401 8415
rect 8435 8381 8447 8415
rect 8389 8375 8447 8381
rect 4982 8304 4988 8356
rect 5040 8344 5046 8356
rect 5353 8347 5411 8353
rect 5353 8344 5365 8347
rect 5040 8316 5365 8344
rect 5040 8304 5046 8316
rect 5353 8313 5365 8316
rect 5399 8313 5411 8347
rect 5353 8307 5411 8313
rect 5736 8316 6316 8344
rect 5736 8285 5764 8316
rect 6288 8288 6316 8316
rect 6380 8288 6408 8375
rect 8404 8344 8432 8375
rect 9784 8353 9812 8452
rect 9861 8449 9873 8452
rect 9907 8449 9919 8483
rect 9861 8443 9919 8449
rect 10042 8440 10048 8492
rect 10100 8440 10106 8492
rect 7668 8316 8432 8344
rect 4632 8248 4927 8276
rect 5721 8279 5779 8285
rect 5721 8245 5733 8279
rect 5767 8245 5779 8279
rect 5721 8239 5779 8245
rect 5902 8236 5908 8288
rect 5960 8236 5966 8288
rect 6270 8236 6276 8288
rect 6328 8236 6334 8288
rect 6362 8236 6368 8288
rect 6420 8276 6426 8288
rect 7668 8276 7696 8316
rect 6420 8248 7696 8276
rect 8404 8276 8432 8316
rect 9769 8347 9827 8353
rect 9769 8313 9781 8347
rect 9815 8313 9827 8347
rect 9769 8307 9827 8313
rect 8570 8276 8576 8288
rect 8404 8248 8576 8276
rect 6420 8236 6426 8248
rect 8570 8236 8576 8248
rect 8628 8236 8634 8288
rect 1104 8186 12788 8208
rect 1104 8134 2410 8186
rect 2462 8134 2474 8186
rect 2526 8134 2538 8186
rect 2590 8134 2602 8186
rect 2654 8134 2666 8186
rect 2718 8134 5331 8186
rect 5383 8134 5395 8186
rect 5447 8134 5459 8186
rect 5511 8134 5523 8186
rect 5575 8134 5587 8186
rect 5639 8134 8252 8186
rect 8304 8134 8316 8186
rect 8368 8134 8380 8186
rect 8432 8134 8444 8186
rect 8496 8134 8508 8186
rect 8560 8134 11173 8186
rect 11225 8134 11237 8186
rect 11289 8134 11301 8186
rect 11353 8134 11365 8186
rect 11417 8134 11429 8186
rect 11481 8134 12788 8186
rect 1104 8112 12788 8134
rect 2777 8075 2835 8081
rect 2777 8041 2789 8075
rect 2823 8072 2835 8075
rect 3326 8072 3332 8084
rect 2823 8044 3332 8072
rect 2823 8041 2835 8044
rect 2777 8035 2835 8041
rect 3326 8032 3332 8044
rect 3384 8032 3390 8084
rect 3970 8032 3976 8084
rect 4028 8072 4034 8084
rect 4890 8072 4896 8084
rect 4028 8044 4896 8072
rect 4028 8032 4034 8044
rect 4890 8032 4896 8044
rect 4948 8032 4954 8084
rect 10042 8032 10048 8084
rect 10100 8072 10106 8084
rect 10321 8075 10379 8081
rect 10321 8072 10333 8075
rect 10100 8044 10333 8072
rect 10100 8032 10106 8044
rect 10321 8041 10333 8044
rect 10367 8041 10379 8075
rect 10321 8035 10379 8041
rect 1394 7896 1400 7948
rect 1452 7896 1458 7948
rect 5721 7939 5779 7945
rect 5721 7905 5733 7939
rect 5767 7936 5779 7939
rect 7098 7936 7104 7948
rect 5767 7908 7104 7936
rect 5767 7905 5779 7908
rect 5721 7899 5779 7905
rect 7098 7896 7104 7908
rect 7156 7896 7162 7948
rect 8570 7896 8576 7948
rect 8628 7936 8634 7948
rect 8941 7939 8999 7945
rect 8941 7936 8953 7939
rect 8628 7908 8953 7936
rect 8628 7896 8634 7908
rect 8941 7905 8953 7908
rect 8987 7905 8999 7939
rect 8941 7899 8999 7905
rect 1664 7871 1722 7877
rect 1664 7837 1676 7871
rect 1710 7868 1722 7871
rect 2130 7868 2136 7880
rect 1710 7840 2136 7868
rect 1710 7837 1722 7840
rect 1664 7831 1722 7837
rect 2130 7828 2136 7840
rect 2188 7828 2194 7880
rect 3878 7828 3884 7880
rect 3936 7828 3942 7880
rect 4062 7828 4068 7880
rect 4120 7828 4126 7880
rect 4522 7828 4528 7880
rect 4580 7868 4586 7880
rect 4580 7840 4844 7868
rect 4580 7828 4586 7840
rect 4816 7812 4844 7840
rect 5810 7828 5816 7880
rect 5868 7828 5874 7880
rect 7742 7828 7748 7880
rect 7800 7868 7806 7880
rect 7837 7871 7895 7877
rect 7837 7868 7849 7871
rect 7800 7840 7849 7868
rect 7800 7828 7806 7840
rect 7837 7837 7849 7840
rect 7883 7837 7895 7871
rect 7837 7831 7895 7837
rect 8110 7828 8116 7880
rect 8168 7828 8174 7880
rect 3973 7803 4031 7809
rect 3973 7769 3985 7803
rect 4019 7800 4031 7803
rect 4614 7800 4620 7812
rect 4019 7772 4620 7800
rect 4019 7769 4031 7772
rect 3973 7763 4031 7769
rect 4614 7760 4620 7772
rect 4672 7760 4678 7812
rect 4798 7760 4804 7812
rect 4856 7760 4862 7812
rect 6270 7760 6276 7812
rect 6328 7800 6334 7812
rect 7650 7800 7656 7812
rect 6328 7772 7656 7800
rect 6328 7760 6334 7772
rect 7650 7760 7656 7772
rect 7708 7760 7714 7812
rect 9208 7803 9266 7809
rect 9208 7769 9220 7803
rect 9254 7800 9266 7803
rect 9306 7800 9312 7812
rect 9254 7772 9312 7800
rect 9254 7769 9266 7772
rect 9208 7763 9266 7769
rect 9306 7760 9312 7772
rect 9364 7760 9370 7812
rect 4338 7692 4344 7744
rect 4396 7732 4402 7744
rect 4433 7735 4491 7741
rect 4433 7732 4445 7735
rect 4396 7704 4445 7732
rect 4396 7692 4402 7704
rect 4433 7701 4445 7704
rect 4479 7701 4491 7735
rect 4433 7695 4491 7701
rect 5074 7692 5080 7744
rect 5132 7692 5138 7744
rect 5350 7692 5356 7744
rect 5408 7732 5414 7744
rect 7101 7735 7159 7741
rect 7101 7732 7113 7735
rect 5408 7704 7113 7732
rect 5408 7692 5414 7704
rect 7101 7701 7113 7704
rect 7147 7701 7159 7735
rect 7101 7695 7159 7701
rect 1104 7642 12788 7664
rect 1104 7590 3070 7642
rect 3122 7590 3134 7642
rect 3186 7590 3198 7642
rect 3250 7590 3262 7642
rect 3314 7590 3326 7642
rect 3378 7590 5991 7642
rect 6043 7590 6055 7642
rect 6107 7590 6119 7642
rect 6171 7590 6183 7642
rect 6235 7590 6247 7642
rect 6299 7590 8912 7642
rect 8964 7590 8976 7642
rect 9028 7590 9040 7642
rect 9092 7590 9104 7642
rect 9156 7590 9168 7642
rect 9220 7590 11833 7642
rect 11885 7590 11897 7642
rect 11949 7590 11961 7642
rect 12013 7590 12025 7642
rect 12077 7590 12089 7642
rect 12141 7590 12788 7642
rect 1104 7568 12788 7590
rect 1394 7488 1400 7540
rect 1452 7488 1458 7540
rect 4798 7488 4804 7540
rect 4856 7528 4862 7540
rect 5813 7531 5871 7537
rect 5813 7528 5825 7531
rect 4856 7500 5825 7528
rect 4856 7488 4862 7500
rect 5813 7497 5825 7500
rect 5859 7497 5871 7531
rect 5813 7491 5871 7497
rect 5902 7488 5908 7540
rect 5960 7488 5966 7540
rect 7745 7531 7803 7537
rect 7745 7497 7757 7531
rect 7791 7528 7803 7531
rect 7834 7528 7840 7540
rect 7791 7500 7840 7528
rect 7791 7497 7803 7500
rect 7745 7491 7803 7497
rect 7834 7488 7840 7500
rect 7892 7488 7898 7540
rect 10965 7531 11023 7537
rect 10965 7497 10977 7531
rect 11011 7497 11023 7531
rect 10965 7491 11023 7497
rect 1412 7460 1440 7488
rect 2593 7463 2651 7469
rect 2593 7460 2605 7463
rect 1412 7432 2605 7460
rect 2593 7429 2605 7432
rect 2639 7429 2651 7463
rect 2593 7423 2651 7429
rect 4341 7463 4399 7469
rect 4341 7429 4353 7463
rect 4387 7460 4399 7463
rect 5166 7460 5172 7472
rect 4387 7432 5172 7460
rect 4387 7429 4399 7432
rect 4341 7423 4399 7429
rect 5166 7420 5172 7432
rect 5224 7460 5230 7472
rect 5350 7460 5356 7472
rect 5224 7432 5356 7460
rect 5224 7420 5230 7432
rect 5350 7420 5356 7432
rect 5408 7420 5414 7472
rect 4522 7352 4528 7404
rect 4580 7392 4586 7404
rect 4689 7395 4747 7401
rect 4689 7392 4701 7395
rect 4580 7364 4701 7392
rect 4580 7352 4586 7364
rect 4689 7361 4701 7364
rect 4735 7361 4747 7395
rect 4689 7355 4747 7361
rect 4982 7352 4988 7404
rect 5040 7392 5046 7404
rect 5920 7392 5948 7488
rect 6632 7463 6690 7469
rect 6632 7429 6644 7463
rect 6678 7460 6690 7463
rect 7190 7460 7196 7472
rect 6678 7432 7196 7460
rect 6678 7429 6690 7432
rect 6632 7423 6690 7429
rect 7190 7420 7196 7432
rect 7248 7420 7254 7472
rect 9024 7463 9082 7469
rect 7760 7432 8156 7460
rect 7760 7404 7788 7432
rect 5997 7395 6055 7401
rect 5997 7392 6009 7395
rect 5040 7364 5886 7392
rect 5920 7364 6009 7392
rect 5040 7352 5046 7364
rect 4430 7284 4436 7336
rect 4488 7284 4494 7336
rect 5858 7324 5886 7364
rect 5997 7361 6009 7364
rect 6043 7361 6055 7395
rect 5997 7355 6055 7361
rect 6362 7352 6368 7404
rect 6420 7352 6426 7404
rect 6472 7364 7696 7392
rect 6472 7324 6500 7364
rect 5858 7296 6500 7324
rect 7668 7324 7696 7364
rect 7742 7352 7748 7404
rect 7800 7352 7806 7404
rect 7929 7395 7987 7401
rect 7929 7361 7941 7395
rect 7975 7392 7987 7395
rect 8018 7392 8024 7404
rect 7975 7364 8024 7392
rect 7975 7361 7987 7364
rect 7929 7355 7987 7361
rect 8018 7352 8024 7364
rect 8076 7352 8082 7404
rect 8128 7401 8156 7432
rect 9024 7429 9036 7463
rect 9070 7460 9082 7463
rect 10980 7460 11008 7491
rect 9070 7432 11008 7460
rect 9070 7429 9082 7432
rect 9024 7423 9082 7429
rect 8113 7395 8171 7401
rect 8113 7361 8125 7395
rect 8159 7361 8171 7395
rect 8113 7355 8171 7361
rect 8297 7395 8355 7401
rect 8297 7361 8309 7395
rect 8343 7361 8355 7395
rect 8297 7355 8355 7361
rect 8481 7395 8539 7401
rect 8481 7361 8493 7395
rect 8527 7392 8539 7395
rect 8846 7392 8852 7404
rect 8527 7364 8852 7392
rect 8527 7361 8539 7364
rect 8481 7355 8539 7361
rect 8312 7324 8340 7355
rect 8846 7352 8852 7364
rect 8904 7352 8910 7404
rect 9582 7352 9588 7404
rect 9640 7392 9646 7404
rect 10229 7395 10287 7401
rect 10229 7392 10241 7395
rect 9640 7364 10241 7392
rect 9640 7352 9646 7364
rect 10229 7361 10241 7364
rect 10275 7361 10287 7395
rect 10229 7355 10287 7361
rect 11054 7352 11060 7404
rect 11112 7392 11118 7404
rect 11149 7395 11207 7401
rect 11149 7392 11161 7395
rect 11112 7364 11161 7392
rect 11112 7352 11118 7364
rect 11149 7361 11161 7364
rect 11195 7361 11207 7395
rect 11149 7355 11207 7361
rect 8570 7324 8576 7336
rect 7668 7296 8576 7324
rect 8570 7284 8576 7296
rect 8628 7284 8634 7336
rect 8662 7284 8668 7336
rect 8720 7284 8726 7336
rect 8754 7284 8760 7336
rect 8812 7284 8818 7336
rect 10781 7327 10839 7333
rect 10781 7324 10793 7327
rect 10152 7296 10793 7324
rect 2222 7148 2228 7200
rect 2280 7148 2286 7200
rect 2498 7148 2504 7200
rect 2556 7148 2562 7200
rect 6181 7191 6239 7197
rect 6181 7157 6193 7191
rect 6227 7188 6239 7191
rect 7282 7188 7288 7200
rect 6227 7160 7288 7188
rect 6227 7157 6239 7160
rect 6181 7151 6239 7157
rect 7282 7148 7288 7160
rect 7340 7148 7346 7200
rect 9766 7148 9772 7200
rect 9824 7188 9830 7200
rect 10152 7197 10180 7296
rect 10781 7293 10793 7296
rect 10827 7293 10839 7327
rect 10781 7287 10839 7293
rect 10137 7191 10195 7197
rect 10137 7188 10149 7191
rect 9824 7160 10149 7188
rect 9824 7148 9830 7160
rect 10137 7157 10149 7160
rect 10183 7157 10195 7191
rect 10137 7151 10195 7157
rect 1104 7098 12788 7120
rect 1104 7046 2410 7098
rect 2462 7046 2474 7098
rect 2526 7046 2538 7098
rect 2590 7046 2602 7098
rect 2654 7046 2666 7098
rect 2718 7046 5331 7098
rect 5383 7046 5395 7098
rect 5447 7046 5459 7098
rect 5511 7046 5523 7098
rect 5575 7046 5587 7098
rect 5639 7046 8252 7098
rect 8304 7046 8316 7098
rect 8368 7046 8380 7098
rect 8432 7046 8444 7098
rect 8496 7046 8508 7098
rect 8560 7046 11173 7098
rect 11225 7046 11237 7098
rect 11289 7046 11301 7098
rect 11353 7046 11365 7098
rect 11417 7046 11429 7098
rect 11481 7046 12788 7098
rect 1104 7024 12788 7046
rect 3605 6987 3663 6993
rect 3605 6953 3617 6987
rect 3651 6984 3663 6987
rect 3881 6987 3939 6993
rect 3881 6984 3893 6987
rect 3651 6956 3893 6984
rect 3651 6953 3663 6956
rect 3605 6947 3663 6953
rect 3881 6953 3893 6956
rect 3927 6984 3939 6987
rect 4062 6984 4068 6996
rect 3927 6956 4068 6984
rect 3927 6953 3939 6956
rect 3881 6947 3939 6953
rect 4062 6944 4068 6956
rect 4120 6944 4126 6996
rect 6362 6944 6368 6996
rect 6420 6984 6426 6996
rect 6549 6987 6607 6993
rect 6549 6984 6561 6987
rect 6420 6956 6561 6984
rect 6420 6944 6426 6956
rect 6549 6953 6561 6956
rect 6595 6953 6607 6987
rect 6549 6947 6607 6953
rect 8662 6944 8668 6996
rect 8720 6984 8726 6996
rect 8720 6956 9352 6984
rect 8720 6944 8726 6956
rect 3694 6876 3700 6928
rect 3752 6916 3758 6928
rect 4890 6916 4896 6928
rect 3752 6888 4896 6916
rect 3752 6876 3758 6888
rect 4890 6876 4896 6888
rect 4948 6916 4954 6928
rect 7101 6919 7159 6925
rect 7101 6916 7113 6919
rect 4948 6888 7113 6916
rect 4948 6876 4954 6888
rect 3789 6851 3847 6857
rect 3789 6817 3801 6851
rect 3835 6848 3847 6851
rect 3878 6848 3884 6860
rect 3835 6820 3884 6848
rect 3835 6817 3847 6820
rect 3789 6811 3847 6817
rect 3878 6808 3884 6820
rect 3936 6808 3942 6860
rect 3970 6808 3976 6860
rect 4028 6808 4034 6860
rect 4246 6808 4252 6860
rect 4304 6848 4310 6860
rect 4304 6820 5120 6848
rect 4304 6808 4310 6820
rect 1949 6783 2007 6789
rect 1949 6749 1961 6783
rect 1995 6749 2007 6783
rect 1949 6743 2007 6749
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6780 2283 6783
rect 2774 6780 2780 6792
rect 2271 6752 2780 6780
rect 2271 6749 2283 6752
rect 2225 6743 2283 6749
rect 1964 6644 1992 6743
rect 2774 6740 2780 6752
rect 2832 6740 2838 6792
rect 3510 6740 3516 6792
rect 3568 6780 3574 6792
rect 3568 6752 4292 6780
rect 3568 6740 3574 6752
rect 2314 6672 2320 6724
rect 2372 6712 2378 6724
rect 2470 6715 2528 6721
rect 2470 6712 2482 6715
rect 2372 6684 2482 6712
rect 2372 6672 2378 6684
rect 2470 6681 2482 6684
rect 2516 6681 2528 6715
rect 2470 6675 2528 6681
rect 4154 6672 4160 6724
rect 4212 6672 4218 6724
rect 4264 6712 4292 6752
rect 4338 6740 4344 6792
rect 4396 6740 4402 6792
rect 4614 6740 4620 6792
rect 4672 6740 4678 6792
rect 4798 6740 4804 6792
rect 4856 6740 4862 6792
rect 4982 6740 4988 6792
rect 5040 6740 5046 6792
rect 5092 6712 5120 6820
rect 5184 6789 5212 6888
rect 5828 6792 5856 6888
rect 7101 6885 7113 6888
rect 7147 6885 7159 6919
rect 7101 6879 7159 6885
rect 8754 6876 8760 6928
rect 8812 6876 8818 6928
rect 9324 6916 9352 6956
rect 9950 6916 9956 6928
rect 9324 6888 9956 6916
rect 8481 6851 8539 6857
rect 8481 6817 8493 6851
rect 8527 6848 8539 6851
rect 8772 6848 8800 6876
rect 9324 6857 9352 6888
rect 9950 6876 9956 6888
rect 10008 6876 10014 6928
rect 8527 6820 8800 6848
rect 9309 6851 9367 6857
rect 8527 6817 8539 6820
rect 8481 6811 8539 6817
rect 9309 6817 9321 6851
rect 9355 6817 9367 6851
rect 9309 6811 9367 6817
rect 9493 6851 9551 6857
rect 9493 6817 9505 6851
rect 9539 6848 9551 6851
rect 12250 6848 12256 6860
rect 9539 6820 12256 6848
rect 9539 6817 9551 6820
rect 9493 6811 9551 6817
rect 12250 6808 12256 6820
rect 12308 6808 12314 6860
rect 5169 6783 5227 6789
rect 5169 6749 5181 6783
rect 5215 6749 5227 6783
rect 5169 6743 5227 6749
rect 5258 6740 5264 6792
rect 5316 6780 5322 6792
rect 5316 6752 5361 6780
rect 5316 6740 5322 6752
rect 5810 6740 5816 6792
rect 5868 6740 5874 6792
rect 7282 6740 7288 6792
rect 7340 6780 7346 6792
rect 8214 6783 8272 6789
rect 8214 6780 8226 6783
rect 7340 6752 8226 6780
rect 7340 6740 7346 6752
rect 8214 6749 8226 6752
rect 8260 6749 8272 6783
rect 8214 6743 8272 6749
rect 8757 6783 8815 6789
rect 8757 6749 8769 6783
rect 8803 6780 8815 6783
rect 8803 6752 9444 6780
rect 8803 6749 8815 6752
rect 8757 6743 8815 6749
rect 8846 6712 8852 6724
rect 4264 6684 4844 6712
rect 5092 6684 8852 6712
rect 3418 6644 3424 6656
rect 1964 6616 3424 6644
rect 3418 6604 3424 6616
rect 3476 6604 3482 6656
rect 4065 6647 4123 6653
rect 4065 6613 4077 6647
rect 4111 6644 4123 6647
rect 4706 6644 4712 6656
rect 4111 6616 4712 6644
rect 4111 6613 4123 6616
rect 4065 6607 4123 6613
rect 4706 6604 4712 6616
rect 4764 6604 4770 6656
rect 4816 6644 4844 6684
rect 8846 6672 8852 6684
rect 8904 6712 8910 6724
rect 9306 6712 9312 6724
rect 8904 6684 9312 6712
rect 8904 6672 8910 6684
rect 9306 6672 9312 6684
rect 9364 6672 9370 6724
rect 9416 6656 9444 6752
rect 9582 6740 9588 6792
rect 9640 6740 9646 6792
rect 11054 6740 11060 6792
rect 11112 6740 11118 6792
rect 5718 6644 5724 6656
rect 4816 6616 5724 6644
rect 5718 6604 5724 6616
rect 5776 6604 5782 6656
rect 8662 6604 8668 6656
rect 8720 6604 8726 6656
rect 9398 6604 9404 6656
rect 9456 6604 9462 6656
rect 9953 6647 10011 6653
rect 9953 6613 9965 6647
rect 9999 6644 10011 6647
rect 11072 6644 11100 6740
rect 9999 6616 11100 6644
rect 9999 6613 10011 6616
rect 9953 6607 10011 6613
rect 1104 6554 12788 6576
rect 1104 6502 3070 6554
rect 3122 6502 3134 6554
rect 3186 6502 3198 6554
rect 3250 6502 3262 6554
rect 3314 6502 3326 6554
rect 3378 6502 5991 6554
rect 6043 6502 6055 6554
rect 6107 6502 6119 6554
rect 6171 6502 6183 6554
rect 6235 6502 6247 6554
rect 6299 6502 8912 6554
rect 8964 6502 8976 6554
rect 9028 6502 9040 6554
rect 9092 6502 9104 6554
rect 9156 6502 9168 6554
rect 9220 6502 11833 6554
rect 11885 6502 11897 6554
rect 11949 6502 11961 6554
rect 12013 6502 12025 6554
rect 12077 6502 12089 6554
rect 12141 6502 12788 6554
rect 1104 6480 12788 6502
rect 1857 6443 1915 6449
rect 1857 6409 1869 6443
rect 1903 6440 1915 6443
rect 3421 6443 3479 6449
rect 1903 6412 2774 6440
rect 1903 6409 1915 6412
rect 1857 6403 1915 6409
rect 2314 6381 2320 6384
rect 2286 6375 2320 6381
rect 1780 6344 2084 6372
rect 1780 6313 1808 6344
rect 1765 6307 1823 6313
rect 1765 6273 1777 6307
rect 1811 6273 1823 6307
rect 1765 6267 1823 6273
rect 1949 6307 2007 6313
rect 1949 6273 1961 6307
rect 1995 6273 2007 6307
rect 2056 6304 2084 6344
rect 2286 6341 2298 6375
rect 2286 6335 2320 6341
rect 2314 6332 2320 6335
rect 2372 6332 2378 6384
rect 2746 6372 2774 6412
rect 3421 6409 3433 6443
rect 3467 6440 3479 6443
rect 3878 6440 3884 6452
rect 3467 6412 3884 6440
rect 3467 6409 3479 6412
rect 3421 6403 3479 6409
rect 3878 6400 3884 6412
rect 3936 6400 3942 6452
rect 4798 6440 4804 6452
rect 3988 6412 4804 6440
rect 3988 6372 4016 6412
rect 4798 6400 4804 6412
rect 4856 6400 4862 6452
rect 4890 6400 4896 6452
rect 4948 6440 4954 6452
rect 4948 6412 6767 6440
rect 4948 6400 4954 6412
rect 4522 6372 4528 6384
rect 2746 6344 4016 6372
rect 4080 6344 4528 6372
rect 2056 6276 3464 6304
rect 1949 6267 2007 6273
rect 1964 6112 1992 6267
rect 2041 6239 2099 6245
rect 2041 6205 2053 6239
rect 2087 6205 2099 6239
rect 2041 6199 2099 6205
rect 1670 6060 1676 6112
rect 1728 6060 1734 6112
rect 1946 6060 1952 6112
rect 2004 6060 2010 6112
rect 2056 6100 2084 6199
rect 3436 6168 3464 6276
rect 3510 6264 3516 6316
rect 3568 6264 3574 6316
rect 3694 6264 3700 6316
rect 3752 6264 3758 6316
rect 3786 6264 3792 6316
rect 3844 6264 3850 6316
rect 3878 6264 3884 6316
rect 3936 6264 3942 6316
rect 4080 6313 4108 6344
rect 4522 6332 4528 6344
rect 4580 6332 4586 6384
rect 4700 6375 4758 6381
rect 4700 6341 4712 6375
rect 4746 6372 4758 6375
rect 5074 6372 5080 6384
rect 4746 6344 5080 6372
rect 4746 6341 4758 6344
rect 4700 6335 4758 6341
rect 5074 6332 5080 6344
rect 5132 6332 5138 6384
rect 5997 6375 6055 6381
rect 5997 6341 6009 6375
rect 6043 6372 6055 6375
rect 6362 6372 6368 6384
rect 6043 6344 6368 6372
rect 6043 6341 6055 6344
rect 5997 6335 6055 6341
rect 6362 6332 6368 6344
rect 6420 6332 6426 6384
rect 4065 6307 4123 6313
rect 4065 6273 4077 6307
rect 4111 6273 4123 6307
rect 4065 6267 4123 6273
rect 4157 6307 4215 6313
rect 4157 6273 4169 6307
rect 4203 6304 4215 6307
rect 4338 6304 4344 6316
rect 4203 6276 4344 6304
rect 4203 6273 4215 6276
rect 4157 6267 4215 6273
rect 4338 6264 4344 6276
rect 4396 6264 4402 6316
rect 4430 6264 4436 6316
rect 4488 6264 4494 6316
rect 4540 6276 5764 6304
rect 4249 6239 4307 6245
rect 4249 6205 4261 6239
rect 4295 6236 4307 6239
rect 4540 6236 4568 6276
rect 4295 6208 4568 6236
rect 5736 6236 5764 6276
rect 5902 6264 5908 6316
rect 5960 6264 5966 6316
rect 6178 6264 6184 6316
rect 6236 6264 6242 6316
rect 6365 6239 6423 6245
rect 6365 6236 6377 6239
rect 5736 6208 6377 6236
rect 4295 6205 4307 6208
rect 4249 6199 4307 6205
rect 3970 6168 3976 6180
rect 3436 6140 3976 6168
rect 3970 6128 3976 6140
rect 4028 6128 4034 6180
rect 5736 6168 5764 6208
rect 6365 6205 6377 6208
rect 6411 6236 6423 6239
rect 6638 6236 6644 6248
rect 6411 6208 6644 6236
rect 6411 6205 6423 6208
rect 6365 6199 6423 6205
rect 6638 6196 6644 6208
rect 6696 6196 6702 6248
rect 6739 6236 6767 6412
rect 7098 6400 7104 6452
rect 7156 6400 7162 6452
rect 7834 6400 7840 6452
rect 7892 6440 7898 6452
rect 9125 6443 9183 6449
rect 9125 6440 9137 6443
rect 7892 6412 9137 6440
rect 7892 6400 7898 6412
rect 9125 6409 9137 6412
rect 9171 6409 9183 6443
rect 9125 6403 9183 6409
rect 10042 6400 10048 6452
rect 10100 6440 10106 6452
rect 10229 6443 10287 6449
rect 10229 6440 10241 6443
rect 10100 6412 10241 6440
rect 10100 6400 10106 6412
rect 10229 6409 10241 6412
rect 10275 6409 10287 6443
rect 10229 6403 10287 6409
rect 9628 6372 9634 6384
rect 8772 6344 9634 6372
rect 7009 6307 7067 6313
rect 7009 6273 7021 6307
rect 7055 6304 7067 6307
rect 7377 6307 7435 6313
rect 7377 6304 7389 6307
rect 7055 6276 7389 6304
rect 7055 6273 7067 6276
rect 7009 6267 7067 6273
rect 7377 6273 7389 6276
rect 7423 6273 7435 6307
rect 7377 6267 7435 6273
rect 7558 6264 7564 6316
rect 7616 6304 7622 6316
rect 7745 6307 7803 6313
rect 7745 6304 7757 6307
rect 7616 6276 7757 6304
rect 7616 6264 7622 6276
rect 7745 6273 7757 6276
rect 7791 6273 7803 6307
rect 8018 6304 8024 6316
rect 7745 6267 7803 6273
rect 7852 6276 8024 6304
rect 7285 6239 7343 6245
rect 7285 6236 7297 6239
rect 6739 6208 7297 6236
rect 7285 6205 7297 6208
rect 7331 6236 7343 6239
rect 7852 6236 7880 6276
rect 8018 6264 8024 6276
rect 8076 6264 8082 6316
rect 8110 6264 8116 6316
rect 8168 6264 8174 6316
rect 8772 6313 8800 6344
rect 9628 6332 9634 6344
rect 9686 6332 9692 6384
rect 9858 6332 9864 6384
rect 9916 6372 9922 6384
rect 10137 6375 10195 6381
rect 9916 6344 10088 6372
rect 9916 6332 9922 6344
rect 8757 6307 8815 6313
rect 8588 6302 8699 6304
rect 8496 6276 8699 6302
rect 8496 6274 8616 6276
rect 7331 6208 7880 6236
rect 7331 6205 7343 6208
rect 7285 6199 7343 6205
rect 8202 6196 8208 6248
rect 8260 6196 8266 6248
rect 8496 6236 8524 6274
rect 8671 6245 8699 6276
rect 8757 6273 8769 6307
rect 8803 6273 8815 6307
rect 8757 6267 8815 6273
rect 8846 6264 8852 6316
rect 8904 6264 8910 6316
rect 9030 6264 9036 6316
rect 9088 6264 9094 6316
rect 9306 6264 9312 6316
rect 9364 6264 9370 6316
rect 10060 6304 10088 6344
rect 10137 6341 10149 6375
rect 10183 6372 10195 6375
rect 10183 6344 11284 6372
rect 10183 6341 10195 6344
rect 10137 6335 10195 6341
rect 11256 6313 11284 6344
rect 10413 6307 10471 6313
rect 10413 6304 10425 6307
rect 9416 6276 9674 6304
rect 10060 6276 10425 6304
rect 8312 6208 8524 6236
rect 8665 6239 8723 6245
rect 5813 6171 5871 6177
rect 5813 6168 5825 6171
rect 5736 6140 5825 6168
rect 5813 6137 5825 6140
rect 5859 6137 5871 6171
rect 5813 6131 5871 6137
rect 6089 6171 6147 6177
rect 6089 6137 6101 6171
rect 6135 6168 6147 6171
rect 8312 6168 8340 6208
rect 8665 6205 8677 6239
rect 8711 6205 8723 6239
rect 8864 6236 8892 6264
rect 9416 6236 9444 6276
rect 8864 6208 9444 6236
rect 8665 6199 8723 6205
rect 9490 6196 9496 6248
rect 9548 6196 9554 6248
rect 9646 6236 9674 6276
rect 10413 6273 10425 6276
rect 10459 6273 10471 6307
rect 10413 6267 10471 6273
rect 10781 6307 10839 6313
rect 10781 6273 10793 6307
rect 10827 6304 10839 6307
rect 11241 6307 11299 6313
rect 10827 6276 11008 6304
rect 10827 6273 10839 6276
rect 10781 6267 10839 6273
rect 9858 6236 9864 6248
rect 9646 6208 9864 6236
rect 9858 6196 9864 6208
rect 9916 6196 9922 6248
rect 10226 6196 10232 6248
rect 10284 6236 10290 6248
rect 10689 6239 10747 6245
rect 10689 6236 10701 6239
rect 10284 6208 10701 6236
rect 10284 6196 10290 6208
rect 10689 6205 10701 6208
rect 10735 6236 10747 6239
rect 10873 6239 10931 6245
rect 10873 6236 10885 6239
rect 10735 6208 10885 6236
rect 10735 6205 10747 6208
rect 10689 6199 10747 6205
rect 10873 6205 10885 6208
rect 10919 6205 10931 6239
rect 10873 6199 10931 6205
rect 6135 6140 8340 6168
rect 8481 6171 8539 6177
rect 6135 6137 6147 6140
rect 6089 6131 6147 6137
rect 8481 6137 8493 6171
rect 8527 6137 8539 6171
rect 8481 6131 8539 6137
rect 2774 6100 2780 6112
rect 2056 6072 2780 6100
rect 2774 6060 2780 6072
rect 2832 6060 2838 6112
rect 3789 6103 3847 6109
rect 3789 6069 3801 6103
rect 3835 6100 3847 6103
rect 4062 6100 4068 6112
rect 3835 6072 4068 6100
rect 3835 6069 3847 6072
rect 3789 6063 3847 6069
rect 4062 6060 4068 6072
rect 4120 6060 4126 6112
rect 4341 6103 4399 6109
rect 4341 6069 4353 6103
rect 4387 6100 4399 6103
rect 5074 6100 5080 6112
rect 4387 6072 5080 6100
rect 4387 6069 4399 6072
rect 4341 6063 4399 6069
rect 5074 6060 5080 6072
rect 5132 6060 5138 6112
rect 7926 6060 7932 6112
rect 7984 6100 7990 6112
rect 8496 6100 8524 6131
rect 9306 6128 9312 6180
rect 9364 6168 9370 6180
rect 10980 6168 11008 6276
rect 11241 6273 11253 6307
rect 11287 6273 11299 6307
rect 11241 6267 11299 6273
rect 9364 6140 11008 6168
rect 9364 6128 9370 6140
rect 7984 6072 8524 6100
rect 7984 6060 7990 6072
rect 8938 6060 8944 6112
rect 8996 6100 9002 6112
rect 10597 6103 10655 6109
rect 10597 6100 10609 6103
rect 8996 6072 10609 6100
rect 8996 6060 9002 6072
rect 10597 6069 10609 6072
rect 10643 6069 10655 6103
rect 10597 6063 10655 6069
rect 11054 6060 11060 6112
rect 11112 6060 11118 6112
rect 1104 6010 12788 6032
rect 1104 5958 2410 6010
rect 2462 5958 2474 6010
rect 2526 5958 2538 6010
rect 2590 5958 2602 6010
rect 2654 5958 2666 6010
rect 2718 5958 5331 6010
rect 5383 5958 5395 6010
rect 5447 5958 5459 6010
rect 5511 5958 5523 6010
rect 5575 5958 5587 6010
rect 5639 5958 8252 6010
rect 8304 5958 8316 6010
rect 8368 5958 8380 6010
rect 8432 5958 8444 6010
rect 8496 5958 8508 6010
rect 8560 5958 11173 6010
rect 11225 5958 11237 6010
rect 11289 5958 11301 6010
rect 11353 5958 11365 6010
rect 11417 5958 11429 6010
rect 11481 5958 12788 6010
rect 1104 5936 12788 5958
rect 1670 5856 1676 5908
rect 1728 5856 1734 5908
rect 3510 5896 3516 5908
rect 1964 5868 3516 5896
rect 1688 5624 1716 5856
rect 1964 5701 1992 5868
rect 3510 5856 3516 5868
rect 3568 5856 3574 5908
rect 3605 5899 3663 5905
rect 3605 5865 3617 5899
rect 3651 5896 3663 5899
rect 3970 5896 3976 5908
rect 3651 5868 3976 5896
rect 3651 5865 3663 5868
rect 3605 5859 3663 5865
rect 3970 5856 3976 5868
rect 4028 5856 4034 5908
rect 4062 5856 4068 5908
rect 4120 5896 4126 5908
rect 4890 5896 4896 5908
rect 4120 5868 4896 5896
rect 4120 5856 4126 5868
rect 4890 5856 4896 5868
rect 4948 5856 4954 5908
rect 5074 5856 5080 5908
rect 5132 5856 5138 5908
rect 5445 5899 5503 5905
rect 5445 5865 5457 5899
rect 5491 5896 5503 5899
rect 5902 5896 5908 5908
rect 5491 5868 5908 5896
rect 5491 5865 5503 5868
rect 5445 5859 5503 5865
rect 5902 5856 5908 5868
rect 5960 5856 5966 5908
rect 6638 5856 6644 5908
rect 6696 5896 6702 5908
rect 8021 5899 8079 5905
rect 6696 5868 7972 5896
rect 6696 5856 6702 5868
rect 5092 5760 5120 5856
rect 6914 5828 6920 5840
rect 5828 5800 6920 5828
rect 5092 5732 5672 5760
rect 1949 5695 2007 5701
rect 1949 5661 1961 5695
rect 1995 5661 2007 5695
rect 1949 5655 2007 5661
rect 2130 5652 2136 5704
rect 2188 5652 2194 5704
rect 2225 5695 2283 5701
rect 2225 5661 2237 5695
rect 2271 5692 2283 5695
rect 2774 5692 2780 5704
rect 2271 5664 2780 5692
rect 2271 5661 2283 5664
rect 2225 5655 2283 5661
rect 2774 5652 2780 5664
rect 2832 5692 2838 5704
rect 3789 5695 3847 5701
rect 3789 5692 3801 5695
rect 2832 5664 3801 5692
rect 2832 5652 2838 5664
rect 3789 5661 3801 5664
rect 3835 5692 3847 5695
rect 4430 5692 4436 5704
rect 3835 5664 4436 5692
rect 3835 5661 3847 5664
rect 3789 5655 3847 5661
rect 4430 5652 4436 5664
rect 4488 5652 4494 5704
rect 5644 5701 5672 5732
rect 5828 5701 5856 5800
rect 6914 5788 6920 5800
rect 6972 5788 6978 5840
rect 7024 5800 7696 5828
rect 5997 5763 6055 5769
rect 5997 5760 6009 5763
rect 5920 5732 6009 5760
rect 5920 5704 5948 5732
rect 5997 5729 6009 5732
rect 6043 5729 6055 5763
rect 6178 5760 6184 5772
rect 5997 5723 6055 5729
rect 6104 5732 6184 5760
rect 5261 5695 5319 5701
rect 5261 5692 5273 5695
rect 4917 5664 5273 5692
rect 2470 5627 2528 5633
rect 2470 5624 2482 5627
rect 1688 5596 2482 5624
rect 2470 5593 2482 5596
rect 2516 5593 2528 5627
rect 2470 5587 2528 5593
rect 3418 5584 3424 5636
rect 3476 5624 3482 5636
rect 4034 5627 4092 5633
rect 4034 5624 4046 5627
rect 3476 5596 4046 5624
rect 3476 5584 3482 5596
rect 4034 5593 4046 5596
rect 4080 5593 4092 5627
rect 4034 5587 4092 5593
rect 4246 5584 4252 5636
rect 4304 5624 4310 5636
rect 4917 5624 4945 5664
rect 5261 5661 5273 5664
rect 5307 5661 5319 5695
rect 5261 5655 5319 5661
rect 5353 5695 5411 5701
rect 5353 5661 5365 5695
rect 5399 5661 5411 5695
rect 5353 5655 5411 5661
rect 5629 5695 5687 5701
rect 5629 5661 5641 5695
rect 5675 5661 5687 5695
rect 5629 5655 5687 5661
rect 5813 5695 5871 5701
rect 5813 5661 5825 5695
rect 5859 5661 5871 5695
rect 5813 5655 5871 5661
rect 4304 5596 4945 5624
rect 4304 5584 4310 5596
rect 4982 5584 4988 5636
rect 5040 5624 5046 5636
rect 5368 5624 5396 5655
rect 5902 5652 5908 5704
rect 5960 5652 5966 5704
rect 6104 5701 6132 5732
rect 6178 5720 6184 5732
rect 6236 5760 6242 5772
rect 6362 5760 6368 5772
rect 6236 5732 6368 5760
rect 6236 5720 6242 5732
rect 6362 5720 6368 5732
rect 6420 5760 6426 5772
rect 7024 5760 7052 5800
rect 7377 5763 7435 5769
rect 7377 5760 7389 5763
rect 6420 5732 7052 5760
rect 7116 5732 7389 5760
rect 6420 5720 6426 5732
rect 7116 5704 7144 5732
rect 7377 5729 7389 5732
rect 7423 5729 7435 5763
rect 7377 5723 7435 5729
rect 7668 5760 7696 5800
rect 7944 5760 7972 5868
rect 8021 5865 8033 5899
rect 8067 5896 8079 5899
rect 8110 5896 8116 5908
rect 8067 5868 8116 5896
rect 8067 5865 8079 5868
rect 8021 5859 8079 5865
rect 8110 5856 8116 5868
rect 8168 5856 8174 5908
rect 11054 5896 11060 5908
rect 10152 5868 11060 5896
rect 8846 5828 8852 5840
rect 8404 5800 8852 5828
rect 8404 5772 8432 5800
rect 8846 5788 8852 5800
rect 8904 5788 8910 5840
rect 8205 5763 8263 5769
rect 8205 5760 8217 5763
rect 7668 5732 7880 5760
rect 7944 5732 8217 5760
rect 7668 5704 7696 5732
rect 6089 5695 6147 5701
rect 6089 5661 6101 5695
rect 6135 5661 6147 5695
rect 6089 5655 6147 5661
rect 6454 5652 6460 5704
rect 6512 5652 6518 5704
rect 6638 5652 6644 5704
rect 6696 5652 6702 5704
rect 7098 5652 7104 5704
rect 7156 5652 7162 5704
rect 7282 5652 7288 5704
rect 7340 5652 7346 5704
rect 7650 5652 7656 5704
rect 7708 5652 7714 5704
rect 7742 5652 7748 5704
rect 7800 5652 7806 5704
rect 7852 5692 7880 5732
rect 8205 5729 8217 5732
rect 8251 5729 8263 5763
rect 8205 5723 8263 5729
rect 8386 5720 8392 5772
rect 8444 5720 8450 5772
rect 8754 5720 8760 5772
rect 8812 5760 8818 5772
rect 9033 5763 9091 5769
rect 9033 5760 9045 5763
rect 8812 5732 9045 5760
rect 8812 5720 8818 5732
rect 9033 5729 9045 5732
rect 9079 5729 9091 5763
rect 9033 5723 9091 5729
rect 7948 5695 8006 5701
rect 7948 5692 7960 5695
rect 7852 5664 7960 5692
rect 7948 5661 7960 5664
rect 7994 5661 8006 5695
rect 7948 5655 8006 5661
rect 8110 5652 8116 5704
rect 8168 5652 8174 5704
rect 8297 5695 8355 5701
rect 8297 5661 8309 5695
rect 8343 5692 8355 5695
rect 8662 5692 8668 5704
rect 8343 5664 8668 5692
rect 8343 5661 8355 5664
rect 8297 5655 8355 5661
rect 5040 5596 5396 5624
rect 5537 5627 5595 5633
rect 5040 5584 5046 5596
rect 5537 5593 5549 5627
rect 5583 5624 5595 5627
rect 8312 5624 8340 5655
rect 8662 5652 8668 5664
rect 8720 5652 8726 5704
rect 9300 5695 9358 5701
rect 9300 5661 9312 5695
rect 9346 5692 9358 5695
rect 10152 5692 10180 5868
rect 11054 5856 11060 5868
rect 11112 5856 11118 5908
rect 10502 5720 10508 5772
rect 10560 5760 10566 5772
rect 11057 5763 11115 5769
rect 11057 5760 11069 5763
rect 10560 5732 11069 5760
rect 10560 5720 10566 5732
rect 11057 5729 11069 5732
rect 11103 5729 11115 5763
rect 11057 5723 11115 5729
rect 9346 5664 10180 5692
rect 9346 5661 9358 5664
rect 9300 5655 9358 5661
rect 10318 5652 10324 5704
rect 10376 5692 10382 5704
rect 11425 5695 11483 5701
rect 11425 5692 11437 5695
rect 10376 5664 11437 5692
rect 10376 5652 10382 5664
rect 11425 5661 11437 5664
rect 11471 5661 11483 5695
rect 11425 5655 11483 5661
rect 8573 5627 8631 5633
rect 8573 5624 8585 5627
rect 5583 5596 8340 5624
rect 8404 5596 8585 5624
rect 5583 5593 5595 5596
rect 5537 5587 5595 5593
rect 1486 5516 1492 5568
rect 1544 5556 1550 5568
rect 1949 5559 2007 5565
rect 1949 5556 1961 5559
rect 1544 5528 1961 5556
rect 1544 5516 1550 5528
rect 1949 5525 1961 5528
rect 1995 5525 2007 5559
rect 1949 5519 2007 5525
rect 2038 5516 2044 5568
rect 2096 5556 2102 5568
rect 4154 5556 4160 5568
rect 2096 5528 4160 5556
rect 2096 5516 2102 5528
rect 4154 5516 4160 5528
rect 4212 5556 4218 5568
rect 5169 5559 5227 5565
rect 5169 5556 5181 5559
rect 4212 5528 5181 5556
rect 4212 5516 4218 5528
rect 5169 5525 5181 5528
rect 5215 5525 5227 5559
rect 5169 5519 5227 5525
rect 6641 5559 6699 5565
rect 6641 5525 6653 5559
rect 6687 5556 6699 5559
rect 6730 5556 6736 5568
rect 6687 5528 6736 5556
rect 6687 5525 6699 5528
rect 6641 5519 6699 5525
rect 6730 5516 6736 5528
rect 6788 5556 6794 5568
rect 7742 5556 7748 5568
rect 6788 5528 7748 5556
rect 6788 5516 6794 5528
rect 7742 5516 7748 5528
rect 7800 5516 7806 5568
rect 7834 5516 7840 5568
rect 7892 5516 7898 5568
rect 8018 5516 8024 5568
rect 8076 5556 8082 5568
rect 8404 5556 8432 5596
rect 8573 5593 8585 5596
rect 8619 5593 8631 5627
rect 8573 5587 8631 5593
rect 9582 5584 9588 5636
rect 9640 5624 9646 5636
rect 9640 5596 11284 5624
rect 9640 5584 9646 5596
rect 8076 5528 8432 5556
rect 8481 5559 8539 5565
rect 8076 5516 8082 5528
rect 8481 5525 8493 5559
rect 8527 5556 8539 5559
rect 9858 5556 9864 5568
rect 8527 5528 9864 5556
rect 8527 5525 8539 5528
rect 8481 5519 8539 5525
rect 9858 5516 9864 5528
rect 9916 5516 9922 5568
rect 9950 5516 9956 5568
rect 10008 5556 10014 5568
rect 10318 5556 10324 5568
rect 10008 5528 10324 5556
rect 10008 5516 10014 5528
rect 10318 5516 10324 5528
rect 10376 5516 10382 5568
rect 10410 5516 10416 5568
rect 10468 5516 10474 5568
rect 10502 5516 10508 5568
rect 10560 5516 10566 5568
rect 11256 5565 11284 5596
rect 11241 5559 11299 5565
rect 11241 5525 11253 5559
rect 11287 5525 11299 5559
rect 11241 5519 11299 5525
rect 1104 5466 12788 5488
rect 1104 5414 3070 5466
rect 3122 5414 3134 5466
rect 3186 5414 3198 5466
rect 3250 5414 3262 5466
rect 3314 5414 3326 5466
rect 3378 5414 5991 5466
rect 6043 5414 6055 5466
rect 6107 5414 6119 5466
rect 6171 5414 6183 5466
rect 6235 5414 6247 5466
rect 6299 5414 8912 5466
rect 8964 5414 8976 5466
rect 9028 5414 9040 5466
rect 9092 5414 9104 5466
rect 9156 5414 9168 5466
rect 9220 5414 11833 5466
rect 11885 5414 11897 5466
rect 11949 5414 11961 5466
rect 12013 5414 12025 5466
rect 12077 5414 12089 5466
rect 12141 5414 12788 5466
rect 1104 5392 12788 5414
rect 5902 5352 5908 5364
rect 4264 5324 5908 5352
rect 4154 5284 4160 5296
rect 2240 5256 4160 5284
rect 2240 5225 2268 5256
rect 4154 5244 4160 5256
rect 4212 5244 4218 5296
rect 1857 5219 1915 5225
rect 1857 5185 1869 5219
rect 1903 5185 1915 5219
rect 1857 5179 1915 5185
rect 2225 5219 2283 5225
rect 2225 5185 2237 5219
rect 2271 5185 2283 5219
rect 2409 5219 2467 5225
rect 2409 5216 2421 5219
rect 2225 5179 2283 5185
rect 2332 5188 2421 5216
rect 1872 5080 1900 5179
rect 2332 5080 2360 5188
rect 2409 5185 2421 5188
rect 2455 5185 2467 5219
rect 2409 5179 2467 5185
rect 2501 5219 2559 5225
rect 2501 5185 2513 5219
rect 2547 5216 2559 5219
rect 4264 5216 4292 5324
rect 5902 5312 5908 5324
rect 5960 5352 5966 5364
rect 6178 5352 6184 5364
rect 5960 5324 6184 5352
rect 5960 5312 5966 5324
rect 4341 5287 4399 5293
rect 4341 5253 4353 5287
rect 4387 5284 4399 5287
rect 5166 5284 5172 5296
rect 4387 5256 5172 5284
rect 4387 5253 4399 5256
rect 4341 5247 4399 5253
rect 5166 5244 5172 5256
rect 5224 5244 5230 5296
rect 2547 5188 4292 5216
rect 2547 5185 2559 5188
rect 2501 5179 2559 5185
rect 5074 5176 5080 5228
rect 5132 5216 5138 5228
rect 6012 5225 6040 5324
rect 6178 5312 6184 5324
rect 6236 5312 6242 5364
rect 6362 5312 6368 5364
rect 6420 5352 6426 5364
rect 6549 5355 6607 5361
rect 6549 5352 6561 5355
rect 6420 5324 6561 5352
rect 6420 5312 6426 5324
rect 6549 5321 6561 5324
rect 6595 5321 6607 5355
rect 6549 5315 6607 5321
rect 6641 5355 6699 5361
rect 6641 5321 6653 5355
rect 6687 5352 6699 5355
rect 6914 5352 6920 5364
rect 6687 5324 6920 5352
rect 6687 5321 6699 5324
rect 6641 5315 6699 5321
rect 6914 5312 6920 5324
rect 6972 5352 6978 5364
rect 7834 5352 7840 5364
rect 6972 5324 7840 5352
rect 6972 5312 6978 5324
rect 7834 5312 7840 5324
rect 7892 5312 7898 5364
rect 9401 5355 9459 5361
rect 9401 5321 9413 5355
rect 9447 5352 9459 5355
rect 9490 5352 9496 5364
rect 9447 5324 9496 5352
rect 9447 5321 9459 5324
rect 9401 5315 9459 5321
rect 9490 5312 9496 5324
rect 9548 5312 9554 5364
rect 9769 5355 9827 5361
rect 9769 5321 9781 5355
rect 9815 5352 9827 5355
rect 10502 5352 10508 5364
rect 9815 5324 10508 5352
rect 9815 5321 9827 5324
rect 9769 5315 9827 5321
rect 10502 5312 10508 5324
rect 10560 5312 10566 5364
rect 6730 5247 6736 5296
rect 6717 5244 6736 5247
rect 6788 5244 6794 5296
rect 10321 5287 10379 5293
rect 10321 5284 10333 5287
rect 7300 5256 10333 5284
rect 6717 5241 6775 5244
rect 5638 5219 5696 5225
rect 5638 5216 5650 5219
rect 5132 5188 5650 5216
rect 5132 5176 5138 5188
rect 5638 5185 5650 5188
rect 5684 5185 5696 5219
rect 5638 5179 5696 5185
rect 5997 5219 6055 5225
rect 5997 5185 6009 5219
rect 6043 5185 6055 5219
rect 5997 5179 6055 5185
rect 6181 5219 6239 5225
rect 6181 5185 6193 5219
rect 6227 5216 6239 5219
rect 6270 5216 6276 5228
rect 6227 5188 6276 5216
rect 6227 5185 6239 5188
rect 6181 5179 6239 5185
rect 6270 5176 6276 5188
rect 6328 5176 6334 5228
rect 6454 5176 6460 5228
rect 6512 5176 6518 5228
rect 6717 5207 6729 5241
rect 6763 5207 6775 5241
rect 6717 5201 6775 5207
rect 6914 5176 6920 5228
rect 6972 5216 6978 5228
rect 7300 5225 7328 5256
rect 10321 5253 10333 5256
rect 10367 5253 10379 5287
rect 10321 5247 10379 5253
rect 7009 5219 7067 5225
rect 7009 5216 7021 5219
rect 6972 5188 7021 5216
rect 6972 5176 6978 5188
rect 7009 5185 7021 5188
rect 7055 5185 7067 5219
rect 7009 5179 7067 5185
rect 7285 5219 7343 5225
rect 7285 5185 7297 5219
rect 7331 5185 7343 5219
rect 7285 5179 7343 5185
rect 7653 5219 7711 5225
rect 7653 5185 7665 5219
rect 7699 5185 7711 5219
rect 7653 5179 7711 5185
rect 2774 5108 2780 5160
rect 2832 5108 2838 5160
rect 5905 5151 5963 5157
rect 5905 5117 5917 5151
rect 5951 5117 5963 5151
rect 5905 5111 5963 5117
rect 4798 5080 4804 5092
rect 1872 5052 2176 5080
rect 2332 5052 4804 5080
rect 1670 4972 1676 5024
rect 1728 4972 1734 5024
rect 2038 4972 2044 5024
rect 2096 4972 2102 5024
rect 2148 5012 2176 5052
rect 4798 5040 4804 5052
rect 4856 5040 4862 5092
rect 5920 5080 5948 5111
rect 6086 5108 6092 5160
rect 6144 5148 6150 5160
rect 6365 5151 6423 5157
rect 6365 5148 6377 5151
rect 6144 5120 6377 5148
rect 6144 5108 6150 5120
rect 6365 5117 6377 5120
rect 6411 5148 6423 5151
rect 6472 5148 6500 5176
rect 6825 5151 6883 5157
rect 6411 5120 6767 5148
rect 6411 5117 6423 5120
rect 6365 5111 6423 5117
rect 5920 5052 6408 5080
rect 6380 5024 6408 5052
rect 3418 5012 3424 5024
rect 2148 4984 3424 5012
rect 3418 4972 3424 4984
rect 3476 4972 3482 5024
rect 4338 4972 4344 5024
rect 4396 5012 4402 5024
rect 4525 5015 4583 5021
rect 4525 5012 4537 5015
rect 4396 4984 4537 5012
rect 4396 4972 4402 4984
rect 4525 4981 4537 4984
rect 4571 5012 4583 5015
rect 4614 5012 4620 5024
rect 4571 4984 4620 5012
rect 4571 4981 4583 4984
rect 4525 4975 4583 4981
rect 4614 4972 4620 4984
rect 4672 4972 4678 5024
rect 4982 4972 4988 5024
rect 5040 5012 5046 5024
rect 6089 5015 6147 5021
rect 6089 5012 6101 5015
rect 5040 4984 6101 5012
rect 5040 4972 5046 4984
rect 6089 4981 6101 4984
rect 6135 4981 6147 5015
rect 6089 4975 6147 4981
rect 6362 4972 6368 5024
rect 6420 4972 6426 5024
rect 6638 4972 6644 5024
rect 6696 4972 6702 5024
rect 6739 5012 6767 5120
rect 6825 5117 6837 5151
rect 6871 5148 6883 5151
rect 7668 5148 7696 5179
rect 7742 5176 7748 5228
rect 7800 5176 7806 5228
rect 7834 5176 7840 5228
rect 7892 5176 7898 5228
rect 8113 5219 8171 5225
rect 8113 5185 8125 5219
rect 8159 5185 8171 5219
rect 8113 5179 8171 5185
rect 8481 5219 8539 5225
rect 8481 5185 8493 5219
rect 8527 5185 8539 5219
rect 8481 5179 8539 5185
rect 6871 5120 7696 5148
rect 7760 5148 7788 5176
rect 8128 5148 8156 5179
rect 7760 5120 8156 5148
rect 8496 5148 8524 5179
rect 8570 5176 8576 5228
rect 8628 5216 8634 5228
rect 8757 5219 8815 5225
rect 8757 5216 8769 5219
rect 8628 5188 8769 5216
rect 8628 5176 8634 5188
rect 8757 5185 8769 5188
rect 8803 5185 8815 5219
rect 8757 5179 8815 5185
rect 8938 5176 8944 5228
rect 8996 5176 9002 5228
rect 9214 5176 9220 5228
rect 9272 5216 9278 5228
rect 9582 5216 9588 5228
rect 9272 5188 9588 5216
rect 9272 5176 9278 5188
rect 9582 5176 9588 5188
rect 9640 5176 9646 5228
rect 10410 5176 10416 5228
rect 10468 5214 10474 5228
rect 10468 5186 10511 5214
rect 10468 5176 10474 5186
rect 9766 5148 9772 5160
rect 8496 5120 9772 5148
rect 6871 5117 6883 5120
rect 6825 5111 6883 5117
rect 9766 5108 9772 5120
rect 9824 5148 9830 5160
rect 9861 5151 9919 5157
rect 9861 5148 9873 5151
rect 9824 5120 9873 5148
rect 9824 5108 9830 5120
rect 9861 5117 9873 5120
rect 9907 5117 9919 5151
rect 9861 5111 9919 5117
rect 9950 5108 9956 5160
rect 10008 5108 10014 5160
rect 7098 5040 7104 5092
rect 7156 5040 7162 5092
rect 7193 5083 7251 5089
rect 7193 5049 7205 5083
rect 7239 5080 7251 5083
rect 7282 5080 7288 5092
rect 7239 5052 7288 5080
rect 7239 5049 7251 5052
rect 7193 5043 7251 5049
rect 7282 5040 7288 5052
rect 7340 5080 7346 5092
rect 8573 5083 8631 5089
rect 8573 5080 8585 5083
rect 7340 5052 8585 5080
rect 7340 5040 7346 5052
rect 8573 5049 8585 5052
rect 8619 5049 8631 5083
rect 8573 5043 8631 5049
rect 7466 5012 7472 5024
rect 6739 4984 7472 5012
rect 7466 4972 7472 4984
rect 7524 4972 7530 5024
rect 7742 4972 7748 5024
rect 7800 4972 7806 5024
rect 8386 4972 8392 5024
rect 8444 5012 8450 5024
rect 9490 5012 9496 5024
rect 8444 4984 9496 5012
rect 8444 4972 8450 4984
rect 9490 4972 9496 4984
rect 9548 4972 9554 5024
rect 1104 4922 12788 4944
rect 1104 4870 2410 4922
rect 2462 4870 2474 4922
rect 2526 4870 2538 4922
rect 2590 4870 2602 4922
rect 2654 4870 2666 4922
rect 2718 4870 5331 4922
rect 5383 4870 5395 4922
rect 5447 4870 5459 4922
rect 5511 4870 5523 4922
rect 5575 4870 5587 4922
rect 5639 4870 8252 4922
rect 8304 4870 8316 4922
rect 8368 4870 8380 4922
rect 8432 4870 8444 4922
rect 8496 4870 8508 4922
rect 8560 4870 11173 4922
rect 11225 4870 11237 4922
rect 11289 4870 11301 4922
rect 11353 4870 11365 4922
rect 11417 4870 11429 4922
rect 11481 4870 12788 4922
rect 1104 4848 12788 4870
rect 2038 4768 2044 4820
rect 2096 4808 2102 4820
rect 4709 4811 4767 4817
rect 2096 4780 4476 4808
rect 2096 4768 2102 4780
rect 3510 4700 3516 4752
rect 3568 4740 3574 4752
rect 3786 4740 3792 4752
rect 3568 4712 3792 4740
rect 3568 4700 3574 4712
rect 3786 4700 3792 4712
rect 3844 4700 3850 4752
rect 2590 4632 2596 4684
rect 2648 4672 2654 4684
rect 2961 4675 3019 4681
rect 2961 4672 2973 4675
rect 2648 4644 2973 4672
rect 2648 4632 2654 4644
rect 2961 4641 2973 4644
rect 3007 4641 3019 4675
rect 2961 4635 3019 4641
rect 1397 4607 1455 4613
rect 1397 4573 1409 4607
rect 1443 4604 1455 4607
rect 2774 4604 2780 4616
rect 1443 4576 2780 4604
rect 1443 4573 1455 4576
rect 1397 4567 1455 4573
rect 2774 4564 2780 4576
rect 2832 4564 2838 4616
rect 3605 4607 3663 4613
rect 3605 4573 3617 4607
rect 3651 4604 3663 4607
rect 3694 4604 3700 4616
rect 3651 4576 3700 4604
rect 3651 4573 3663 4576
rect 3605 4567 3663 4573
rect 3694 4564 3700 4576
rect 3752 4564 3758 4616
rect 4338 4564 4344 4616
rect 4396 4564 4402 4616
rect 4448 4604 4476 4780
rect 4709 4777 4721 4811
rect 4755 4808 4767 4811
rect 5442 4808 5448 4820
rect 4755 4780 5448 4808
rect 4755 4777 4767 4780
rect 4709 4771 4767 4777
rect 5442 4768 5448 4780
rect 5500 4768 5506 4820
rect 5718 4808 5724 4820
rect 5644 4780 5724 4808
rect 4893 4743 4951 4749
rect 4893 4709 4905 4743
rect 4939 4740 4951 4743
rect 4939 4712 5488 4740
rect 4939 4709 4951 4712
rect 4893 4703 4951 4709
rect 4985 4675 5043 4681
rect 4985 4641 4997 4675
rect 5031 4672 5043 4675
rect 5074 4672 5080 4684
rect 5031 4644 5080 4672
rect 5031 4641 5043 4644
rect 4985 4635 5043 4641
rect 5074 4632 5080 4644
rect 5132 4632 5138 4684
rect 5460 4681 5488 4712
rect 5445 4675 5503 4681
rect 5445 4641 5457 4675
rect 5491 4641 5503 4675
rect 5445 4635 5503 4641
rect 5534 4632 5540 4684
rect 5592 4632 5598 4684
rect 5169 4607 5227 4613
rect 5169 4604 5181 4607
rect 4448 4576 5181 4604
rect 5169 4573 5181 4576
rect 5215 4573 5227 4607
rect 5169 4567 5227 4573
rect 5258 4564 5264 4616
rect 5316 4564 5322 4616
rect 5353 4607 5411 4613
rect 5353 4573 5365 4607
rect 5399 4604 5411 4607
rect 5552 4604 5580 4632
rect 5644 4613 5672 4780
rect 5718 4768 5724 4780
rect 5776 4768 5782 4820
rect 6454 4808 6460 4820
rect 6104 4780 6460 4808
rect 5810 4632 5816 4684
rect 5868 4672 5874 4684
rect 5997 4675 6055 4681
rect 5997 4672 6009 4675
rect 5868 4644 6009 4672
rect 5868 4632 5874 4644
rect 5997 4641 6009 4644
rect 6043 4641 6055 4675
rect 5997 4635 6055 4641
rect 5399 4576 5580 4604
rect 5629 4607 5687 4613
rect 5399 4573 5411 4576
rect 5353 4567 5411 4573
rect 5629 4573 5641 4607
rect 5675 4573 5687 4607
rect 5629 4567 5687 4573
rect 5721 4607 5779 4613
rect 5721 4573 5733 4607
rect 5767 4604 5779 4607
rect 6104 4604 6132 4780
rect 6454 4768 6460 4780
rect 6512 4768 6518 4820
rect 7004 4780 8984 4808
rect 7004 4740 7032 4780
rect 8956 4752 8984 4780
rect 9306 4768 9312 4820
rect 9364 4768 9370 4820
rect 9490 4768 9496 4820
rect 9548 4768 9554 4820
rect 9766 4768 9772 4820
rect 9824 4768 9830 4820
rect 9858 4768 9864 4820
rect 9916 4768 9922 4820
rect 6380 4712 7032 4740
rect 5767 4576 6132 4604
rect 5767 4573 5779 4576
rect 5721 4567 5779 4573
rect 6178 4564 6184 4616
rect 6236 4564 6242 4616
rect 6270 4564 6276 4616
rect 6328 4564 6334 4616
rect 1670 4545 1676 4548
rect 1664 4536 1676 4545
rect 1631 4508 1676 4536
rect 1664 4499 1676 4508
rect 1670 4496 1676 4499
rect 1728 4496 1734 4548
rect 2038 4496 2044 4548
rect 2096 4536 2102 4548
rect 4525 4539 4583 4545
rect 2096 4508 2912 4536
rect 2096 4496 2102 4508
rect 1946 4428 1952 4480
rect 2004 4468 2010 4480
rect 2130 4468 2136 4480
rect 2004 4440 2136 4468
rect 2004 4428 2010 4440
rect 2130 4428 2136 4440
rect 2188 4468 2194 4480
rect 2682 4468 2688 4480
rect 2188 4440 2688 4468
rect 2188 4428 2194 4440
rect 2682 4428 2688 4440
rect 2740 4468 2746 4480
rect 2777 4471 2835 4477
rect 2777 4468 2789 4471
rect 2740 4440 2789 4468
rect 2740 4428 2746 4440
rect 2777 4437 2789 4440
rect 2823 4437 2835 4471
rect 2884 4468 2912 4508
rect 4525 4505 4537 4539
rect 4571 4536 4583 4539
rect 5534 4536 5540 4548
rect 4571 4508 5540 4536
rect 4571 4505 4583 4508
rect 4525 4499 4583 4505
rect 5534 4496 5540 4508
rect 5592 4496 5598 4548
rect 6380 4536 6408 4712
rect 6638 4672 6644 4684
rect 6564 4644 6644 4672
rect 6564 4613 6592 4644
rect 6638 4632 6644 4644
rect 6696 4632 6702 4684
rect 6549 4607 6607 4613
rect 6549 4573 6561 4607
rect 6595 4573 6607 4607
rect 6549 4567 6607 4573
rect 6917 4607 6975 4613
rect 6917 4573 6929 4607
rect 6963 4604 6975 4607
rect 7004 4604 7032 4712
rect 8110 4700 8116 4752
rect 8168 4700 8174 4752
rect 8938 4700 8944 4752
rect 8996 4700 9002 4752
rect 9324 4740 9352 4768
rect 9140 4712 9352 4740
rect 8021 4675 8079 4681
rect 8021 4641 8033 4675
rect 8067 4672 8079 4675
rect 8128 4672 8156 4700
rect 9140 4681 9168 4712
rect 9125 4675 9183 4681
rect 9125 4672 9137 4675
rect 8067 4644 8156 4672
rect 8772 4644 9137 4672
rect 8067 4641 8079 4644
rect 8021 4635 8079 4641
rect 6963 4576 7032 4604
rect 6963 4573 6975 4576
rect 6917 4567 6975 4573
rect 7466 4564 7472 4616
rect 7524 4564 7530 4616
rect 7650 4564 7656 4616
rect 7708 4604 7714 4616
rect 7745 4607 7803 4613
rect 7745 4604 7757 4607
rect 7708 4576 7757 4604
rect 7708 4564 7714 4576
rect 7745 4573 7757 4576
rect 7791 4573 7803 4607
rect 7745 4567 7803 4573
rect 7834 4564 7840 4616
rect 7892 4604 7898 4616
rect 8113 4607 8171 4613
rect 8113 4604 8125 4607
rect 7892 4576 8125 4604
rect 7892 4564 7898 4576
rect 8113 4573 8125 4576
rect 8159 4573 8171 4607
rect 8113 4567 8171 4573
rect 8478 4564 8484 4616
rect 8536 4564 8542 4616
rect 8772 4613 8800 4644
rect 9125 4641 9137 4644
rect 9171 4641 9183 4675
rect 9125 4635 9183 4641
rect 9214 4632 9220 4684
rect 9272 4632 9278 4684
rect 8757 4607 8815 4613
rect 8757 4573 8769 4607
rect 8803 4573 8815 4607
rect 8757 4567 8815 4573
rect 9300 4607 9358 4613
rect 9300 4573 9312 4607
rect 9346 4573 9358 4607
rect 9300 4567 9358 4573
rect 9401 4607 9459 4613
rect 9401 4573 9413 4607
rect 9447 4604 9459 4607
rect 9508 4604 9536 4768
rect 9674 4632 9680 4684
rect 9732 4672 9738 4684
rect 9769 4675 9827 4681
rect 9769 4672 9781 4675
rect 9732 4644 9781 4672
rect 9732 4632 9738 4644
rect 9769 4641 9781 4644
rect 9815 4641 9827 4675
rect 9769 4635 9827 4641
rect 9447 4576 9536 4604
rect 9953 4607 10011 4613
rect 9447 4573 9459 4576
rect 9401 4567 9459 4573
rect 9953 4573 9965 4607
rect 9999 4604 10011 4607
rect 10042 4604 10048 4616
rect 9999 4576 10048 4604
rect 9999 4573 10011 4576
rect 9953 4567 10011 4573
rect 5644 4508 6408 4536
rect 6457 4539 6515 4545
rect 4614 4468 4620 4480
rect 2884 4440 4620 4468
rect 2777 4431 2835 4437
rect 4614 4428 4620 4440
rect 4672 4468 4678 4480
rect 4735 4471 4793 4477
rect 4735 4468 4747 4471
rect 4672 4440 4747 4468
rect 4672 4428 4678 4440
rect 4735 4437 4747 4440
rect 4781 4468 4793 4471
rect 5350 4468 5356 4480
rect 4781 4440 5356 4468
rect 4781 4437 4793 4440
rect 4735 4431 4793 4437
rect 5350 4428 5356 4440
rect 5408 4468 5414 4480
rect 5644 4468 5672 4508
rect 6457 4505 6469 4539
rect 6503 4536 6515 4539
rect 6822 4536 6828 4548
rect 6503 4508 6828 4536
rect 6503 4505 6515 4508
rect 6457 4499 6515 4505
rect 6822 4496 6828 4508
rect 6880 4496 6886 4548
rect 7484 4536 7512 4564
rect 8018 4536 8024 4548
rect 7484 4508 8024 4536
rect 8018 4496 8024 4508
rect 8076 4536 8082 4548
rect 8496 4536 8524 4564
rect 9315 4536 9343 4567
rect 10042 4564 10048 4576
rect 10100 4564 10106 4616
rect 10226 4564 10232 4616
rect 10284 4564 10290 4616
rect 8076 4508 9343 4536
rect 8076 4496 8082 4508
rect 5408 4440 5672 4468
rect 5813 4471 5871 4477
rect 5408 4428 5414 4440
rect 5813 4437 5825 4471
rect 5859 4468 5871 4471
rect 5902 4468 5908 4480
rect 5859 4440 5908 4468
rect 5859 4437 5871 4440
rect 5813 4431 5871 4437
rect 5902 4428 5908 4440
rect 5960 4428 5966 4480
rect 5997 4471 6055 4477
rect 5997 4437 6009 4471
rect 6043 4468 6055 4471
rect 7558 4468 7564 4480
rect 6043 4440 7564 4468
rect 6043 4437 6055 4440
rect 5997 4431 6055 4437
rect 7558 4428 7564 4440
rect 7616 4428 7622 4480
rect 8662 4428 8668 4480
rect 8720 4468 8726 4480
rect 8941 4471 8999 4477
rect 8941 4468 8953 4471
rect 8720 4440 8953 4468
rect 8720 4428 8726 4440
rect 8941 4437 8953 4440
rect 8987 4437 8999 4471
rect 9315 4468 9343 4508
rect 9582 4496 9588 4548
rect 9640 4496 9646 4548
rect 9398 4468 9404 4480
rect 9315 4440 9404 4468
rect 8941 4431 8999 4437
rect 9398 4428 9404 4440
rect 9456 4428 9462 4480
rect 10042 4428 10048 4480
rect 10100 4428 10106 4480
rect 1104 4378 12788 4400
rect 1104 4326 3070 4378
rect 3122 4326 3134 4378
rect 3186 4326 3198 4378
rect 3250 4326 3262 4378
rect 3314 4326 3326 4378
rect 3378 4326 5991 4378
rect 6043 4326 6055 4378
rect 6107 4326 6119 4378
rect 6171 4326 6183 4378
rect 6235 4326 6247 4378
rect 6299 4326 8912 4378
rect 8964 4326 8976 4378
rect 9028 4326 9040 4378
rect 9092 4326 9104 4378
rect 9156 4326 9168 4378
rect 9220 4326 11833 4378
rect 11885 4326 11897 4378
rect 11949 4326 11961 4378
rect 12013 4326 12025 4378
rect 12077 4326 12089 4378
rect 12141 4326 12788 4378
rect 1104 4304 12788 4326
rect 2774 4224 2780 4276
rect 2832 4264 2838 4276
rect 3053 4267 3111 4273
rect 2832 4236 2912 4264
rect 2832 4224 2838 4236
rect 2590 4156 2596 4208
rect 2648 4196 2654 4208
rect 2694 4199 2752 4205
rect 2694 4196 2706 4199
rect 2648 4168 2706 4196
rect 2648 4156 2654 4168
rect 2694 4165 2706 4168
rect 2740 4165 2752 4199
rect 2694 4159 2752 4165
rect 2884 4128 2912 4236
rect 3053 4233 3065 4267
rect 3099 4264 3111 4267
rect 3418 4264 3424 4276
rect 3099 4236 3424 4264
rect 3099 4233 3111 4236
rect 3053 4227 3111 4233
rect 3418 4224 3424 4236
rect 3476 4224 3482 4276
rect 3602 4224 3608 4276
rect 3660 4264 3666 4276
rect 3881 4267 3939 4273
rect 3881 4264 3893 4267
rect 3660 4236 3893 4264
rect 3660 4224 3666 4236
rect 3881 4233 3893 4236
rect 3927 4233 3939 4267
rect 4614 4264 4620 4276
rect 3881 4227 3939 4233
rect 4060 4236 4620 4264
rect 3142 4156 3148 4208
rect 3200 4196 3206 4208
rect 3237 4199 3295 4205
rect 3237 4196 3249 4199
rect 3200 4168 3249 4196
rect 3200 4156 3206 4168
rect 3237 4165 3249 4168
rect 3283 4165 3295 4199
rect 3237 4159 3295 4165
rect 3697 4199 3755 4205
rect 3697 4165 3709 4199
rect 3743 4196 3755 4199
rect 3786 4196 3792 4208
rect 3743 4168 3792 4196
rect 3743 4165 3755 4168
rect 3697 4159 3755 4165
rect 3786 4156 3792 4168
rect 3844 4156 3850 4208
rect 4060 4137 4088 4236
rect 4614 4224 4620 4236
rect 4672 4224 4678 4276
rect 4982 4224 4988 4276
rect 5040 4224 5046 4276
rect 5077 4267 5135 4273
rect 5077 4233 5089 4267
rect 5123 4264 5135 4267
rect 5258 4264 5264 4276
rect 5123 4236 5264 4264
rect 5123 4233 5135 4236
rect 5077 4227 5135 4233
rect 5258 4224 5264 4236
rect 5316 4224 5322 4276
rect 5350 4224 5356 4276
rect 5408 4264 5414 4276
rect 5445 4267 5503 4273
rect 5445 4264 5457 4267
rect 5408 4236 5457 4264
rect 5408 4224 5414 4236
rect 5445 4233 5457 4236
rect 5491 4233 5503 4267
rect 5445 4227 5503 4233
rect 5534 4224 5540 4276
rect 5592 4264 5598 4276
rect 7742 4264 7748 4276
rect 5592 4236 7748 4264
rect 5592 4224 5598 4236
rect 5000 4196 5028 4224
rect 4172 4168 4476 4196
rect 4172 4140 4200 4168
rect 2961 4131 3019 4137
rect 2961 4128 2973 4131
rect 2884 4100 2973 4128
rect 2961 4097 2973 4100
rect 3007 4097 3019 4131
rect 3957 4131 4015 4137
rect 3957 4128 3969 4131
rect 2961 4091 3019 4097
rect 3896 4100 3969 4128
rect 3605 4063 3663 4069
rect 3605 4029 3617 4063
rect 3651 4060 3663 4063
rect 3896 4060 3924 4100
rect 3957 4097 3969 4100
rect 4003 4097 4015 4131
rect 4060 4131 4123 4137
rect 4060 4100 4077 4131
rect 3957 4091 4015 4097
rect 4065 4097 4077 4100
rect 4111 4097 4123 4131
rect 4065 4091 4123 4097
rect 4154 4088 4160 4140
rect 4212 4088 4218 4140
rect 4448 4137 4476 4168
rect 4724 4168 5212 4196
rect 4724 4137 4752 4168
rect 4249 4131 4307 4137
rect 4249 4097 4261 4131
rect 4295 4097 4307 4131
rect 4249 4091 4307 4097
rect 4341 4131 4399 4137
rect 4341 4097 4353 4131
rect 4387 4097 4399 4131
rect 4341 4091 4399 4097
rect 4433 4131 4491 4137
rect 4433 4097 4445 4131
rect 4479 4097 4491 4131
rect 4433 4091 4491 4097
rect 4709 4131 4767 4137
rect 4709 4097 4721 4131
rect 4755 4097 4767 4131
rect 4709 4091 4767 4097
rect 4801 4131 4859 4137
rect 4801 4097 4813 4131
rect 4847 4128 4859 4131
rect 4890 4128 4896 4140
rect 4847 4100 4896 4128
rect 4847 4097 4859 4100
rect 4801 4091 4859 4097
rect 3651 4032 3924 4060
rect 3651 4029 3663 4032
rect 3605 4023 3663 4029
rect 3694 3952 3700 4004
rect 3752 3952 3758 4004
rect 3896 3992 3924 4032
rect 4264 3992 4292 4091
rect 4356 4060 4384 4091
rect 4890 4088 4896 4100
rect 4948 4088 4954 4140
rect 4985 4131 5043 4137
rect 4985 4097 4997 4131
rect 5031 4128 5043 4131
rect 5074 4128 5080 4140
rect 5031 4100 5080 4128
rect 5031 4097 5043 4100
rect 4985 4091 5043 4097
rect 5074 4088 5080 4100
rect 5132 4088 5138 4140
rect 5184 4128 5212 4168
rect 5261 4131 5319 4137
rect 5261 4128 5273 4131
rect 5184 4100 5273 4128
rect 5261 4097 5273 4100
rect 5307 4097 5319 4131
rect 5261 4091 5319 4097
rect 5442 4088 5448 4140
rect 5500 4128 5506 4140
rect 5537 4131 5595 4137
rect 5537 4128 5549 4131
rect 5500 4100 5549 4128
rect 5500 4088 5506 4100
rect 5537 4097 5549 4100
rect 5583 4097 5595 4131
rect 5537 4091 5595 4097
rect 5552 4060 5580 4091
rect 5626 4088 5632 4140
rect 5684 4088 5690 4140
rect 5736 4128 5764 4236
rect 7742 4224 7748 4236
rect 7800 4224 7806 4276
rect 8938 4264 8944 4276
rect 7852 4236 8944 4264
rect 5813 4199 5871 4205
rect 5813 4165 5825 4199
rect 5859 4196 5871 4199
rect 6822 4196 6828 4208
rect 5859 4168 6828 4196
rect 5859 4165 5871 4168
rect 5813 4159 5871 4165
rect 6822 4156 6828 4168
rect 6880 4156 6886 4208
rect 7098 4156 7104 4208
rect 7156 4196 7162 4208
rect 7852 4196 7880 4236
rect 8938 4224 8944 4236
rect 8996 4224 9002 4276
rect 9033 4267 9091 4273
rect 9033 4233 9045 4267
rect 9079 4264 9091 4267
rect 9490 4264 9496 4276
rect 9079 4236 9496 4264
rect 9079 4233 9091 4236
rect 9033 4227 9091 4233
rect 9490 4224 9496 4236
rect 9548 4224 9554 4276
rect 7156 4168 7880 4196
rect 7156 4156 7162 4168
rect 7926 4156 7932 4208
rect 7984 4196 7990 4208
rect 7984 4168 8248 4196
rect 7984 4156 7990 4168
rect 5905 4131 5963 4137
rect 5905 4128 5917 4131
rect 5736 4100 5917 4128
rect 5905 4097 5917 4100
rect 5951 4097 5963 4131
rect 5905 4091 5963 4097
rect 5997 4131 6055 4137
rect 5997 4097 6009 4131
rect 6043 4128 6055 4131
rect 6043 4100 6132 4128
rect 6043 4097 6055 4100
rect 5997 4091 6055 4097
rect 6104 4060 6132 4100
rect 6454 4088 6460 4140
rect 6512 4128 6518 4140
rect 6621 4131 6679 4137
rect 6621 4128 6633 4131
rect 6512 4100 6633 4128
rect 6512 4088 6518 4100
rect 6621 4097 6633 4100
rect 6667 4097 6679 4131
rect 6840 4128 6868 4156
rect 8220 4137 8248 4168
rect 8478 4156 8484 4208
rect 8536 4196 8542 4208
rect 8536 4168 9076 4196
rect 8536 4156 8542 4168
rect 8113 4131 8171 4137
rect 8113 4128 8125 4131
rect 6840 4100 8125 4128
rect 6621 4091 6679 4097
rect 8113 4097 8125 4100
rect 8159 4097 8171 4131
rect 8113 4091 8171 4097
rect 8205 4131 8263 4137
rect 8205 4097 8217 4131
rect 8251 4097 8263 4131
rect 8205 4091 8263 4097
rect 8573 4131 8631 4137
rect 8573 4097 8585 4131
rect 8619 4097 8631 4131
rect 8573 4091 8631 4097
rect 4356 4032 5488 4060
rect 5552 4032 6132 4060
rect 3896 3964 4200 3992
rect 4264 3964 5120 3992
rect 1581 3927 1639 3933
rect 1581 3893 1593 3927
rect 1627 3924 1639 3927
rect 2222 3924 2228 3936
rect 1627 3896 2228 3924
rect 1627 3893 1639 3896
rect 1581 3887 1639 3893
rect 2222 3884 2228 3896
rect 2280 3884 2286 3936
rect 3237 3927 3295 3933
rect 3237 3893 3249 3927
rect 3283 3924 3295 3927
rect 4062 3924 4068 3936
rect 3283 3896 4068 3924
rect 3283 3893 3295 3896
rect 3237 3887 3295 3893
rect 4062 3884 4068 3896
rect 4120 3884 4126 3936
rect 4172 3924 4200 3964
rect 5092 3936 5120 3964
rect 4246 3924 4252 3936
rect 4172 3896 4252 3924
rect 4246 3884 4252 3896
rect 4304 3884 4310 3936
rect 4614 3884 4620 3936
rect 4672 3884 4678 3936
rect 4982 3884 4988 3936
rect 5040 3884 5046 3936
rect 5074 3884 5080 3936
rect 5132 3884 5138 3936
rect 5460 3924 5488 4032
rect 6104 3936 6132 4032
rect 6362 4020 6368 4072
rect 6420 4020 6426 4072
rect 8588 4060 8616 4091
rect 8662 4088 8668 4140
rect 8720 4088 8726 4140
rect 8772 4137 8800 4168
rect 9048 4140 9076 4168
rect 9306 4156 9312 4208
rect 9364 4156 9370 4208
rect 10042 4156 10048 4208
rect 10100 4156 10106 4208
rect 8757 4131 8815 4137
rect 8757 4097 8769 4131
rect 8803 4097 8815 4131
rect 8757 4091 8815 4097
rect 8846 4088 8852 4140
rect 8904 4088 8910 4140
rect 9030 4088 9036 4140
rect 9088 4088 9094 4140
rect 9125 4131 9183 4137
rect 9125 4097 9137 4131
rect 9171 4128 9183 4131
rect 9324 4128 9352 4156
rect 9171 4100 9352 4128
rect 9484 4131 9542 4137
rect 9171 4097 9183 4100
rect 9125 4091 9183 4097
rect 9484 4097 9496 4131
rect 9530 4128 9542 4131
rect 10060 4128 10088 4156
rect 9530 4100 10088 4128
rect 9530 4097 9542 4100
rect 9484 4091 9542 4097
rect 8864 4060 8892 4088
rect 9217 4063 9275 4069
rect 9217 4060 9229 4063
rect 8588 4032 8708 4060
rect 8864 4032 9229 4060
rect 5718 3924 5724 3936
rect 5460 3896 5724 3924
rect 5718 3884 5724 3896
rect 5776 3884 5782 3936
rect 6086 3884 6092 3936
rect 6144 3884 6150 3936
rect 6181 3927 6239 3933
rect 6181 3893 6193 3927
rect 6227 3924 6239 3927
rect 6270 3924 6276 3936
rect 6227 3896 6276 3924
rect 6227 3893 6239 3896
rect 6181 3887 6239 3893
rect 6270 3884 6276 3896
rect 6328 3884 6334 3936
rect 6380 3924 6408 4020
rect 8680 3992 8708 4032
rect 9217 4029 9229 4032
rect 9263 4029 9275 4063
rect 9217 4023 9275 4029
rect 8849 3995 8907 4001
rect 8849 3992 8861 3995
rect 8680 3964 8861 3992
rect 8849 3961 8861 3964
rect 8895 3961 8907 3995
rect 8849 3955 8907 3961
rect 6730 3924 6736 3936
rect 6380 3896 6736 3924
rect 6730 3884 6736 3896
rect 6788 3884 6794 3936
rect 7006 3884 7012 3936
rect 7064 3924 7070 3936
rect 7650 3924 7656 3936
rect 7064 3896 7656 3924
rect 7064 3884 7070 3896
rect 7650 3884 7656 3896
rect 7708 3924 7714 3936
rect 7745 3927 7803 3933
rect 7745 3924 7757 3927
rect 7708 3896 7757 3924
rect 7708 3884 7714 3896
rect 7745 3893 7757 3896
rect 7791 3893 7803 3927
rect 7745 3887 7803 3893
rect 8297 3927 8355 3933
rect 8297 3893 8309 3927
rect 8343 3924 8355 3927
rect 8662 3924 8668 3936
rect 8343 3896 8668 3924
rect 8343 3893 8355 3896
rect 8297 3887 8355 3893
rect 8662 3884 8668 3896
rect 8720 3884 8726 3936
rect 10594 3884 10600 3936
rect 10652 3884 10658 3936
rect 1104 3834 12788 3856
rect 1104 3782 2410 3834
rect 2462 3782 2474 3834
rect 2526 3782 2538 3834
rect 2590 3782 2602 3834
rect 2654 3782 2666 3834
rect 2718 3782 5331 3834
rect 5383 3782 5395 3834
rect 5447 3782 5459 3834
rect 5511 3782 5523 3834
rect 5575 3782 5587 3834
rect 5639 3782 8252 3834
rect 8304 3782 8316 3834
rect 8368 3782 8380 3834
rect 8432 3782 8444 3834
rect 8496 3782 8508 3834
rect 8560 3782 11173 3834
rect 11225 3782 11237 3834
rect 11289 3782 11301 3834
rect 11353 3782 11365 3834
rect 11417 3782 11429 3834
rect 11481 3782 12788 3834
rect 1104 3760 12788 3782
rect 2130 3680 2136 3732
rect 2188 3720 2194 3732
rect 2188 3692 4200 3720
rect 2188 3680 2194 3692
rect 1397 3655 1455 3661
rect 1397 3621 1409 3655
rect 1443 3652 1455 3655
rect 1443 3624 1808 3652
rect 1443 3621 1455 3624
rect 1397 3615 1455 3621
rect 1780 3516 1808 3624
rect 2777 3587 2835 3593
rect 2777 3553 2789 3587
rect 2823 3584 2835 3587
rect 2866 3584 2872 3596
rect 2823 3556 2872 3584
rect 2823 3553 2835 3556
rect 2777 3547 2835 3553
rect 2866 3544 2872 3556
rect 2924 3544 2930 3596
rect 4172 3593 4200 3692
rect 4614 3680 4620 3732
rect 4672 3680 4678 3732
rect 5718 3680 5724 3732
rect 5776 3720 5782 3732
rect 6546 3720 6552 3732
rect 5776 3692 6552 3720
rect 5776 3680 5782 3692
rect 6546 3680 6552 3692
rect 6604 3680 6610 3732
rect 7101 3723 7159 3729
rect 7101 3689 7113 3723
rect 7147 3689 7159 3723
rect 7101 3683 7159 3689
rect 4157 3587 4215 3593
rect 3344 3556 4016 3584
rect 2682 3516 2688 3528
rect 1780 3488 2688 3516
rect 2682 3476 2688 3488
rect 2740 3516 2746 3528
rect 3344 3516 3372 3556
rect 2740 3488 3372 3516
rect 2740 3476 2746 3488
rect 3418 3476 3424 3528
rect 3476 3476 3482 3528
rect 3988 3525 4016 3556
rect 4157 3553 4169 3587
rect 4203 3584 4215 3587
rect 4338 3584 4344 3596
rect 4203 3556 4344 3584
rect 4203 3553 4215 3556
rect 4157 3547 4215 3553
rect 4338 3544 4344 3556
rect 4396 3544 4402 3596
rect 3973 3519 4031 3525
rect 3973 3485 3985 3519
rect 4019 3485 4031 3519
rect 3973 3479 4031 3485
rect 4065 3519 4123 3525
rect 4065 3485 4077 3519
rect 4111 3485 4123 3519
rect 4065 3479 4123 3485
rect 2532 3451 2590 3457
rect 2532 3417 2544 3451
rect 2578 3448 2590 3451
rect 2869 3451 2927 3457
rect 2869 3448 2881 3451
rect 2578 3420 2881 3448
rect 2578 3417 2590 3420
rect 2532 3411 2590 3417
rect 2869 3417 2881 3420
rect 2915 3417 2927 3451
rect 2869 3411 2927 3417
rect 2958 3408 2964 3460
rect 3016 3448 3022 3460
rect 4080 3448 4108 3479
rect 4246 3476 4252 3528
rect 4304 3476 4310 3528
rect 4433 3519 4491 3525
rect 4433 3485 4445 3519
rect 4479 3516 4491 3519
rect 4632 3516 4660 3680
rect 5902 3612 5908 3664
rect 5960 3652 5966 3664
rect 7116 3652 7144 3683
rect 7282 3680 7288 3732
rect 7340 3720 7346 3732
rect 7742 3720 7748 3732
rect 7340 3692 7748 3720
rect 7340 3680 7346 3692
rect 7742 3680 7748 3692
rect 7800 3720 7806 3732
rect 9033 3723 9091 3729
rect 9033 3720 9045 3723
rect 7800 3692 9045 3720
rect 7800 3680 7806 3692
rect 9033 3689 9045 3692
rect 9079 3689 9091 3723
rect 9033 3683 9091 3689
rect 9401 3723 9459 3729
rect 9401 3689 9413 3723
rect 9447 3720 9459 3723
rect 9582 3720 9588 3732
rect 9447 3692 9588 3720
rect 9447 3689 9459 3692
rect 9401 3683 9459 3689
rect 9582 3680 9588 3692
rect 9640 3680 9646 3732
rect 10226 3680 10232 3732
rect 10284 3720 10290 3732
rect 10413 3723 10471 3729
rect 10413 3720 10425 3723
rect 10284 3692 10425 3720
rect 10284 3680 10290 3692
rect 10413 3689 10425 3692
rect 10459 3689 10471 3723
rect 10413 3683 10471 3689
rect 5960 3624 7144 3652
rect 5960 3612 5966 3624
rect 7466 3612 7472 3664
rect 7524 3652 7530 3664
rect 8110 3652 8116 3664
rect 7524 3624 8116 3652
rect 7524 3612 7530 3624
rect 8110 3612 8116 3624
rect 8168 3652 8174 3664
rect 8168 3624 9260 3652
rect 8168 3612 8174 3624
rect 6730 3544 6736 3596
rect 6788 3584 6794 3596
rect 7009 3587 7067 3593
rect 7009 3584 7021 3587
rect 6788 3556 7021 3584
rect 6788 3544 6794 3556
rect 7009 3553 7021 3556
rect 7055 3584 7067 3587
rect 8754 3584 8760 3596
rect 7055 3556 8760 3584
rect 7055 3553 7067 3556
rect 7009 3547 7067 3553
rect 8754 3544 8760 3556
rect 8812 3544 8818 3596
rect 4479 3488 4660 3516
rect 4479 3485 4491 3488
rect 4433 3479 4491 3485
rect 4706 3476 4712 3528
rect 4764 3476 4770 3528
rect 4798 3476 4804 3528
rect 4856 3525 4862 3528
rect 4856 3519 4883 3525
rect 4871 3485 4883 3519
rect 4856 3479 4883 3485
rect 4856 3476 4862 3479
rect 5166 3476 5172 3528
rect 5224 3516 5230 3528
rect 5261 3519 5319 3525
rect 5261 3516 5273 3519
rect 5224 3488 5273 3516
rect 5224 3476 5230 3488
rect 5261 3485 5273 3488
rect 5307 3485 5319 3519
rect 5261 3479 5319 3485
rect 6086 3476 6092 3528
rect 6144 3516 6150 3528
rect 7466 3516 7472 3528
rect 6144 3488 7472 3516
rect 6144 3476 6150 3488
rect 7466 3476 7472 3488
rect 7524 3476 7530 3528
rect 7650 3476 7656 3528
rect 7708 3476 7714 3528
rect 7926 3476 7932 3528
rect 7984 3516 7990 3528
rect 8481 3519 8539 3525
rect 8481 3516 8493 3519
rect 7984 3488 8493 3516
rect 7984 3476 7990 3488
rect 8481 3485 8493 3488
rect 8527 3516 8539 3519
rect 8570 3516 8576 3528
rect 8527 3488 8576 3516
rect 8527 3485 8539 3488
rect 8481 3479 8539 3485
rect 8570 3476 8576 3488
rect 8628 3516 8634 3528
rect 9232 3525 9260 3624
rect 9490 3544 9496 3596
rect 9548 3584 9554 3596
rect 9769 3587 9827 3593
rect 9769 3584 9781 3587
rect 9548 3556 9781 3584
rect 9548 3544 9554 3556
rect 9769 3553 9781 3556
rect 9815 3553 9827 3587
rect 9769 3547 9827 3553
rect 8941 3519 8999 3525
rect 8941 3516 8953 3519
rect 8628 3488 8953 3516
rect 8628 3476 8634 3488
rect 8941 3485 8953 3488
rect 8987 3485 8999 3519
rect 8941 3479 8999 3485
rect 9217 3519 9275 3525
rect 9217 3485 9229 3519
rect 9263 3516 9275 3519
rect 9306 3516 9312 3528
rect 9263 3488 9312 3516
rect 9263 3485 9275 3488
rect 9217 3479 9275 3485
rect 9306 3476 9312 3488
rect 9364 3476 9370 3528
rect 9953 3519 10011 3525
rect 9953 3485 9965 3519
rect 9999 3516 10011 3519
rect 12250 3516 12256 3528
rect 9999 3488 12256 3516
rect 9999 3485 10011 3488
rect 9953 3479 10011 3485
rect 12250 3476 12256 3488
rect 12308 3476 12314 3528
rect 3016 3420 4568 3448
rect 3016 3408 3022 3420
rect 2314 3340 2320 3392
rect 2372 3380 2378 3392
rect 3789 3383 3847 3389
rect 3789 3380 3801 3383
rect 2372 3352 3801 3380
rect 2372 3340 2378 3352
rect 3789 3349 3801 3352
rect 3835 3349 3847 3383
rect 4540 3380 4568 3420
rect 4614 3408 4620 3460
rect 4672 3408 4678 3460
rect 5718 3448 5724 3460
rect 4917 3420 5724 3448
rect 4917 3380 4945 3420
rect 5718 3408 5724 3420
rect 5776 3408 5782 3460
rect 9030 3408 9036 3460
rect 9088 3448 9094 3460
rect 10045 3451 10103 3457
rect 10045 3448 10057 3451
rect 9088 3420 10057 3448
rect 9088 3408 9094 3420
rect 10045 3417 10057 3420
rect 10091 3448 10103 3451
rect 10594 3448 10600 3460
rect 10091 3420 10600 3448
rect 10091 3417 10103 3420
rect 10045 3411 10103 3417
rect 10594 3408 10600 3420
rect 10652 3408 10658 3460
rect 4540 3352 4945 3380
rect 3789 3343 3847 3349
rect 4982 3340 4988 3392
rect 5040 3340 5046 3392
rect 7926 3340 7932 3392
rect 7984 3340 7990 3392
rect 8938 3340 8944 3392
rect 8996 3380 9002 3392
rect 9490 3380 9496 3392
rect 8996 3352 9496 3380
rect 8996 3340 9002 3352
rect 9490 3340 9496 3352
rect 9548 3340 9554 3392
rect 1104 3290 12788 3312
rect 1104 3238 3070 3290
rect 3122 3238 3134 3290
rect 3186 3238 3198 3290
rect 3250 3238 3262 3290
rect 3314 3238 3326 3290
rect 3378 3238 5991 3290
rect 6043 3238 6055 3290
rect 6107 3238 6119 3290
rect 6171 3238 6183 3290
rect 6235 3238 6247 3290
rect 6299 3238 8912 3290
rect 8964 3238 8976 3290
rect 9028 3238 9040 3290
rect 9092 3238 9104 3290
rect 9156 3238 9168 3290
rect 9220 3238 11833 3290
rect 11885 3238 11897 3290
rect 11949 3238 11961 3290
rect 12013 3238 12025 3290
rect 12077 3238 12089 3290
rect 12141 3238 12788 3290
rect 1104 3216 12788 3238
rect 1857 3179 1915 3185
rect 1857 3145 1869 3179
rect 1903 3176 1915 3179
rect 4522 3176 4528 3188
rect 1903 3148 4528 3176
rect 1903 3145 1915 3148
rect 1857 3139 1915 3145
rect 4522 3136 4528 3148
rect 4580 3136 4586 3188
rect 5074 3176 5080 3188
rect 4632 3148 5080 3176
rect 1578 3068 1584 3120
rect 1636 3068 1642 3120
rect 1765 3111 1823 3117
rect 1765 3077 1777 3111
rect 1811 3108 1823 3111
rect 2314 3108 2320 3120
rect 1811 3080 2320 3108
rect 1811 3077 1823 3080
rect 1765 3071 1823 3077
rect 2314 3068 2320 3080
rect 2372 3068 2378 3120
rect 4632 3108 4660 3148
rect 5074 3136 5080 3148
rect 5132 3176 5138 3188
rect 6089 3179 6147 3185
rect 6089 3176 6101 3179
rect 5132 3148 6101 3176
rect 5132 3136 5138 3148
rect 6089 3145 6101 3148
rect 6135 3145 6147 3179
rect 6089 3139 6147 3145
rect 6362 3136 6368 3188
rect 6420 3136 6426 3188
rect 6457 3179 6515 3185
rect 6457 3145 6469 3179
rect 6503 3176 6515 3179
rect 6546 3176 6552 3188
rect 6503 3148 6552 3176
rect 6503 3145 6515 3148
rect 6457 3139 6515 3145
rect 6546 3136 6552 3148
rect 6604 3136 6610 3188
rect 6638 3136 6644 3188
rect 6696 3176 6702 3188
rect 7653 3179 7711 3185
rect 7653 3176 7665 3179
rect 6696 3148 7665 3176
rect 6696 3136 6702 3148
rect 7653 3145 7665 3148
rect 7699 3145 7711 3179
rect 7653 3139 7711 3145
rect 7926 3136 7932 3188
rect 7984 3136 7990 3188
rect 9401 3179 9459 3185
rect 9401 3145 9413 3179
rect 9447 3176 9459 3179
rect 9490 3176 9496 3188
rect 9447 3148 9496 3176
rect 9447 3145 9459 3148
rect 9401 3139 9459 3145
rect 9490 3136 9496 3148
rect 9548 3136 9554 3188
rect 4798 3108 4804 3120
rect 2608 3080 4660 3108
rect 4724 3080 4804 3108
rect 1486 3000 1492 3052
rect 1544 3000 1550 3052
rect 2038 3000 2044 3052
rect 2096 3000 2102 3052
rect 2225 3043 2283 3049
rect 2225 3009 2237 3043
rect 2271 3040 2283 3043
rect 2608 3040 2636 3080
rect 2271 3012 2636 3040
rect 2271 3009 2283 3012
rect 2225 3003 2283 3009
rect 2682 3000 2688 3052
rect 2740 3000 2746 3052
rect 3050 3000 3056 3052
rect 3108 3000 3114 3052
rect 3418 3000 3424 3052
rect 3476 3000 3482 3052
rect 4246 3040 4252 3052
rect 3712 3012 4252 3040
rect 2130 2932 2136 2984
rect 2188 2972 2194 2984
rect 2317 2975 2375 2981
rect 2317 2972 2329 2975
rect 2188 2944 2329 2972
rect 2188 2932 2194 2944
rect 2317 2941 2329 2944
rect 2363 2972 2375 2975
rect 2700 2972 2728 3000
rect 3436 2972 3464 3000
rect 3712 2984 3740 3012
rect 4246 3000 4252 3012
rect 4304 3000 4310 3052
rect 4430 3000 4436 3052
rect 4488 3040 4494 3052
rect 4724 3049 4752 3080
rect 4798 3068 4804 3080
rect 4856 3068 4862 3120
rect 4982 3068 4988 3120
rect 5040 3108 5046 3120
rect 5902 3108 5908 3120
rect 5040 3080 5304 3108
rect 5040 3068 5046 3080
rect 4709 3043 4767 3049
rect 4709 3042 4721 3043
rect 4704 3040 4721 3042
rect 4488 3012 4721 3040
rect 4488 3000 4494 3012
rect 4709 3009 4721 3012
rect 4755 3009 4767 3043
rect 4709 3003 4767 3009
rect 5074 3000 5080 3052
rect 5132 3000 5138 3052
rect 5276 3049 5304 3080
rect 5552 3080 5908 3108
rect 5552 3049 5580 3080
rect 5902 3068 5908 3080
rect 5960 3068 5966 3120
rect 6380 3108 6408 3136
rect 7282 3108 7288 3120
rect 6380 3080 6868 3108
rect 5261 3043 5319 3049
rect 5261 3009 5273 3043
rect 5307 3009 5319 3043
rect 5261 3003 5319 3009
rect 5537 3043 5595 3049
rect 5537 3009 5549 3043
rect 5583 3009 5595 3043
rect 5537 3003 5595 3009
rect 5718 3000 5724 3052
rect 5776 3040 5782 3052
rect 5997 3043 6055 3049
rect 5997 3040 6009 3043
rect 5776 3012 6009 3040
rect 5776 3000 5782 3012
rect 5997 3009 6009 3012
rect 6043 3009 6055 3043
rect 5997 3003 6055 3009
rect 6086 3000 6092 3052
rect 6144 3040 6150 3052
rect 6365 3043 6423 3049
rect 6365 3040 6377 3043
rect 6144 3012 6377 3040
rect 6144 3000 6150 3012
rect 6365 3009 6377 3012
rect 6411 3009 6423 3043
rect 6365 3003 6423 3009
rect 6454 3000 6460 3052
rect 6512 3000 6518 3052
rect 6638 3000 6644 3052
rect 6696 3000 6702 3052
rect 2363 2944 2728 2972
rect 2792 2944 3464 2972
rect 2363 2941 2375 2944
rect 2317 2935 2375 2941
rect 1765 2907 1823 2913
rect 1765 2873 1777 2907
rect 1811 2904 1823 2907
rect 2792 2904 2820 2944
rect 3694 2932 3700 2984
rect 3752 2932 3758 2984
rect 3789 2975 3847 2981
rect 3789 2941 3801 2975
rect 3835 2941 3847 2975
rect 3789 2935 3847 2941
rect 1811 2876 2820 2904
rect 1811 2873 1823 2876
rect 1765 2867 1823 2873
rect 2866 2864 2872 2916
rect 2924 2904 2930 2916
rect 3804 2904 3832 2935
rect 4522 2932 4528 2984
rect 4580 2972 4586 2984
rect 4893 2975 4951 2981
rect 4893 2972 4905 2975
rect 4580 2944 4905 2972
rect 4580 2932 4586 2944
rect 4893 2941 4905 2944
rect 4939 2941 4951 2975
rect 4893 2935 4951 2941
rect 4982 2932 4988 2984
rect 5040 2932 5046 2984
rect 5629 2975 5687 2981
rect 5629 2941 5641 2975
rect 5675 2972 5687 2975
rect 5810 2972 5816 2984
rect 5675 2944 5816 2972
rect 5675 2941 5687 2944
rect 5629 2935 5687 2941
rect 5810 2932 5816 2944
rect 5868 2932 5874 2984
rect 5905 2975 5963 2981
rect 5905 2941 5917 2975
rect 5951 2972 5963 2975
rect 6472 2972 6500 3000
rect 6840 2981 6868 3080
rect 7208 3080 7288 3108
rect 7208 3049 7236 3080
rect 7282 3068 7288 3080
rect 7340 3068 7346 3120
rect 7466 3068 7472 3120
rect 7524 3068 7530 3120
rect 7944 3108 7972 3136
rect 7760 3080 7972 3108
rect 7193 3043 7251 3049
rect 7193 3009 7205 3043
rect 7239 3009 7251 3043
rect 7193 3003 7251 3009
rect 7377 3043 7435 3049
rect 7377 3009 7389 3043
rect 7423 3040 7435 3043
rect 7484 3040 7512 3068
rect 7760 3049 7788 3080
rect 7423 3012 7512 3040
rect 7745 3043 7803 3049
rect 7423 3009 7435 3012
rect 7377 3003 7435 3009
rect 7745 3009 7757 3043
rect 7791 3009 7803 3043
rect 7745 3003 7803 3009
rect 7837 3043 7895 3049
rect 7837 3009 7849 3043
rect 7883 3040 7895 3043
rect 8754 3040 8760 3052
rect 7883 3012 8760 3040
rect 7883 3009 7895 3012
rect 7837 3003 7895 3009
rect 8754 3000 8760 3012
rect 8812 3000 8818 3052
rect 5951 2944 6500 2972
rect 6825 2975 6883 2981
rect 5951 2941 5963 2944
rect 5905 2935 5963 2941
rect 6825 2941 6837 2975
rect 6871 2941 6883 2975
rect 7285 2975 7343 2981
rect 7285 2972 7297 2975
rect 6825 2935 6883 2941
rect 6932 2944 7297 2972
rect 5994 2904 6000 2916
rect 2924 2876 3832 2904
rect 4356 2876 6000 2904
rect 2924 2864 2930 2876
rect 2961 2839 3019 2845
rect 2961 2805 2973 2839
rect 3007 2836 3019 2839
rect 4356 2836 4384 2876
rect 5994 2864 6000 2876
rect 6052 2864 6058 2916
rect 6733 2907 6791 2913
rect 6733 2873 6745 2907
rect 6779 2904 6791 2907
rect 6932 2904 6960 2944
rect 7285 2941 7297 2944
rect 7331 2941 7343 2975
rect 7285 2935 7343 2941
rect 8113 2975 8171 2981
rect 8113 2941 8125 2975
rect 8159 2972 8171 2975
rect 8570 2972 8576 2984
rect 8159 2944 8576 2972
rect 8159 2941 8171 2944
rect 8113 2935 8171 2941
rect 8570 2932 8576 2944
rect 8628 2932 8634 2984
rect 6779 2876 6960 2904
rect 6779 2873 6791 2876
rect 6733 2867 6791 2873
rect 3007 2808 4384 2836
rect 3007 2805 3019 2808
rect 2961 2799 3019 2805
rect 4430 2796 4436 2848
rect 4488 2796 4494 2848
rect 4522 2796 4528 2848
rect 4580 2796 4586 2848
rect 5810 2796 5816 2848
rect 5868 2836 5874 2848
rect 6748 2836 6776 2867
rect 7006 2864 7012 2916
rect 7064 2864 7070 2916
rect 9674 2904 9680 2916
rect 8772 2876 9680 2904
rect 5868 2808 6776 2836
rect 6825 2839 6883 2845
rect 5868 2796 5874 2808
rect 6825 2805 6837 2839
rect 6871 2836 6883 2839
rect 6914 2836 6920 2848
rect 6871 2808 6920 2836
rect 6871 2805 6883 2808
rect 6825 2799 6883 2805
rect 6914 2796 6920 2808
rect 6972 2796 6978 2848
rect 7024 2836 7052 2864
rect 8772 2836 8800 2876
rect 9674 2864 9680 2876
rect 9732 2864 9738 2916
rect 7024 2808 8800 2836
rect 1104 2746 12788 2768
rect 1104 2694 2410 2746
rect 2462 2694 2474 2746
rect 2526 2694 2538 2746
rect 2590 2694 2602 2746
rect 2654 2694 2666 2746
rect 2718 2694 5331 2746
rect 5383 2694 5395 2746
rect 5447 2694 5459 2746
rect 5511 2694 5523 2746
rect 5575 2694 5587 2746
rect 5639 2694 8252 2746
rect 8304 2694 8316 2746
rect 8368 2694 8380 2746
rect 8432 2694 8444 2746
rect 8496 2694 8508 2746
rect 8560 2694 11173 2746
rect 11225 2694 11237 2746
rect 11289 2694 11301 2746
rect 11353 2694 11365 2746
rect 11417 2694 11429 2746
rect 11481 2694 12788 2746
rect 1104 2672 12788 2694
rect 1946 2592 1952 2644
rect 2004 2632 2010 2644
rect 2133 2635 2191 2641
rect 2133 2632 2145 2635
rect 2004 2604 2145 2632
rect 2004 2592 2010 2604
rect 2133 2601 2145 2604
rect 2179 2601 2191 2635
rect 2133 2595 2191 2601
rect 2777 2635 2835 2641
rect 2777 2601 2789 2635
rect 2823 2632 2835 2635
rect 2866 2632 2872 2644
rect 2823 2604 2872 2632
rect 2823 2601 2835 2604
rect 2777 2595 2835 2601
rect 2866 2592 2872 2604
rect 2924 2592 2930 2644
rect 4522 2632 4528 2644
rect 3344 2604 4528 2632
rect 2222 2456 2228 2508
rect 2280 2456 2286 2508
rect 2314 2456 2320 2508
rect 2372 2496 2378 2508
rect 2593 2499 2651 2505
rect 2593 2496 2605 2499
rect 2372 2468 2605 2496
rect 2372 2456 2378 2468
rect 2593 2465 2605 2468
rect 2639 2465 2651 2499
rect 2593 2459 2651 2465
rect 2130 2388 2136 2440
rect 2188 2437 2194 2440
rect 2188 2428 2196 2437
rect 2188 2400 2233 2428
rect 2188 2391 2196 2400
rect 2188 2388 2194 2391
rect 3050 2388 3056 2440
rect 3108 2388 3114 2440
rect 3344 2437 3372 2604
rect 4522 2592 4528 2604
rect 4580 2592 4586 2644
rect 4798 2592 4804 2644
rect 4856 2632 4862 2644
rect 6457 2635 6515 2641
rect 6457 2632 6469 2635
rect 4856 2604 6469 2632
rect 4856 2592 4862 2604
rect 6457 2601 6469 2604
rect 6503 2601 6515 2635
rect 6457 2595 6515 2601
rect 8110 2592 8116 2644
rect 8168 2592 8174 2644
rect 8570 2592 8576 2644
rect 8628 2592 8634 2644
rect 8662 2592 8668 2644
rect 8720 2592 8726 2644
rect 9030 2592 9036 2644
rect 9088 2592 9094 2644
rect 12250 2592 12256 2644
rect 12308 2592 12314 2644
rect 5442 2524 5448 2576
rect 5500 2564 5506 2576
rect 6086 2564 6092 2576
rect 5500 2536 6092 2564
rect 5500 2524 5506 2536
rect 6086 2524 6092 2536
rect 6144 2524 6150 2576
rect 5169 2499 5227 2505
rect 5169 2465 5181 2499
rect 5215 2496 5227 2499
rect 6730 2496 6736 2508
rect 5215 2468 6736 2496
rect 5215 2465 5227 2468
rect 5169 2459 5227 2465
rect 6730 2456 6736 2468
rect 6788 2456 6794 2508
rect 8481 2499 8539 2505
rect 8481 2465 8493 2499
rect 8527 2465 8539 2499
rect 9398 2496 9404 2508
rect 8481 2459 8539 2465
rect 9048 2468 9404 2496
rect 3329 2431 3387 2437
rect 3329 2397 3341 2431
rect 3375 2397 3387 2431
rect 3329 2391 3387 2397
rect 3605 2431 3663 2437
rect 3605 2397 3617 2431
rect 3651 2428 3663 2431
rect 3878 2428 3884 2440
rect 3651 2400 3884 2428
rect 3651 2397 3663 2400
rect 3605 2391 3663 2397
rect 3878 2388 3884 2400
rect 3936 2428 3942 2440
rect 4154 2428 4160 2440
rect 3936 2400 4160 2428
rect 3936 2388 3942 2400
rect 4154 2388 4160 2400
rect 4212 2388 4218 2440
rect 4430 2388 4436 2440
rect 4488 2428 4494 2440
rect 4902 2431 4960 2437
rect 4902 2428 4914 2431
rect 4488 2400 4914 2428
rect 4488 2388 4494 2400
rect 4902 2397 4914 2400
rect 4948 2397 4960 2431
rect 4902 2391 4960 2397
rect 5629 2431 5687 2437
rect 5629 2397 5641 2431
rect 5675 2428 5687 2431
rect 5718 2428 5724 2440
rect 5675 2400 5724 2428
rect 5675 2397 5687 2400
rect 5629 2391 5687 2397
rect 5718 2388 5724 2400
rect 5776 2388 5782 2440
rect 5810 2388 5816 2440
rect 5868 2388 5874 2440
rect 5994 2388 6000 2440
rect 6052 2428 6058 2440
rect 7006 2437 7012 2440
rect 6365 2431 6423 2437
rect 6365 2428 6377 2431
rect 6052 2400 6377 2428
rect 6052 2388 6058 2400
rect 6365 2397 6377 2400
rect 6411 2397 6423 2431
rect 6365 2391 6423 2397
rect 6989 2431 7012 2437
rect 6989 2397 7001 2431
rect 6989 2391 7012 2397
rect 7006 2388 7012 2391
rect 7064 2388 7070 2440
rect 14 2320 20 2372
rect 72 2360 78 2372
rect 1397 2363 1455 2369
rect 1397 2360 1409 2363
rect 72 2332 1409 2360
rect 72 2320 78 2332
rect 1397 2329 1409 2332
rect 1443 2329 1455 2363
rect 1397 2323 1455 2329
rect 1765 2363 1823 2369
rect 1765 2329 1777 2363
rect 1811 2360 1823 2363
rect 3145 2363 3203 2369
rect 3145 2360 3157 2363
rect 1811 2332 3157 2360
rect 1811 2329 1823 2332
rect 1765 2323 1823 2329
rect 3145 2329 3157 2332
rect 3191 2329 3203 2363
rect 3145 2323 3203 2329
rect 3513 2363 3571 2369
rect 3513 2329 3525 2363
rect 3559 2360 3571 2363
rect 4982 2360 4988 2372
rect 3559 2332 4988 2360
rect 3559 2329 3571 2332
rect 3513 2323 3571 2329
rect 4982 2320 4988 2332
rect 5040 2360 5046 2372
rect 5040 2332 5396 2360
rect 5040 2320 5046 2332
rect 2501 2295 2559 2301
rect 2501 2261 2513 2295
rect 2547 2292 2559 2295
rect 2961 2295 3019 2301
rect 2961 2292 2973 2295
rect 2547 2264 2973 2292
rect 2547 2261 2559 2264
rect 2501 2255 2559 2261
rect 2961 2261 2973 2264
rect 3007 2292 3019 2295
rect 3602 2292 3608 2304
rect 3007 2264 3608 2292
rect 3007 2261 3019 2264
rect 2961 2255 3019 2261
rect 3602 2252 3608 2264
rect 3660 2252 3666 2304
rect 3786 2252 3792 2304
rect 3844 2252 3850 2304
rect 4062 2252 4068 2304
rect 4120 2292 4126 2304
rect 5261 2295 5319 2301
rect 5261 2292 5273 2295
rect 4120 2264 5273 2292
rect 4120 2252 4126 2264
rect 5261 2261 5273 2264
rect 5307 2261 5319 2295
rect 5368 2292 5396 2332
rect 5442 2320 5448 2372
rect 5500 2320 5506 2372
rect 5905 2295 5963 2301
rect 5905 2292 5917 2295
rect 5368 2264 5917 2292
rect 5261 2255 5319 2261
rect 5905 2261 5917 2264
rect 5951 2261 5963 2295
rect 8496 2292 8524 2459
rect 8757 2431 8815 2437
rect 8757 2397 8769 2431
rect 8803 2397 8815 2431
rect 8757 2391 8815 2397
rect 8941 2431 8999 2437
rect 8941 2397 8953 2431
rect 8987 2428 8999 2431
rect 9048 2428 9076 2468
rect 9398 2456 9404 2468
rect 9456 2456 9462 2508
rect 8987 2400 9076 2428
rect 9125 2431 9183 2437
rect 8987 2397 8999 2400
rect 8941 2391 8999 2397
rect 9125 2397 9137 2431
rect 9171 2428 9183 2431
rect 9306 2428 9312 2440
rect 9171 2400 9312 2428
rect 9171 2397 9183 2400
rect 9125 2391 9183 2397
rect 8772 2360 8800 2391
rect 9306 2388 9312 2400
rect 9364 2388 9370 2440
rect 9582 2388 9588 2440
rect 9640 2388 9646 2440
rect 12437 2431 12495 2437
rect 12437 2397 12449 2431
rect 12483 2428 12495 2431
rect 12483 2400 12848 2428
rect 12483 2397 12495 2400
rect 12437 2391 12495 2397
rect 9600 2360 9628 2388
rect 8772 2332 9628 2360
rect 12820 2304 12848 2400
rect 9766 2292 9772 2304
rect 8496 2264 9772 2292
rect 5905 2255 5963 2261
rect 9766 2252 9772 2264
rect 9824 2252 9830 2304
rect 12802 2252 12808 2304
rect 12860 2252 12866 2304
rect 1104 2202 12788 2224
rect 1104 2150 3070 2202
rect 3122 2150 3134 2202
rect 3186 2150 3198 2202
rect 3250 2150 3262 2202
rect 3314 2150 3326 2202
rect 3378 2150 5991 2202
rect 6043 2150 6055 2202
rect 6107 2150 6119 2202
rect 6171 2150 6183 2202
rect 6235 2150 6247 2202
rect 6299 2150 8912 2202
rect 8964 2150 8976 2202
rect 9028 2150 9040 2202
rect 9092 2150 9104 2202
rect 9156 2150 9168 2202
rect 9220 2150 11833 2202
rect 11885 2150 11897 2202
rect 11949 2150 11961 2202
rect 12013 2150 12025 2202
rect 12077 2150 12089 2202
rect 12141 2150 12788 2202
rect 1104 2128 12788 2150
rect 3786 2048 3792 2100
rect 3844 2088 3850 2100
rect 5810 2088 5816 2100
rect 3844 2060 5816 2088
rect 3844 2048 3850 2060
rect 5810 2048 5816 2060
rect 5868 2048 5874 2100
rect 4338 1980 4344 2032
rect 4396 2020 4402 2032
rect 5442 2020 5448 2032
rect 4396 1992 5448 2020
rect 4396 1980 4402 1992
rect 5442 1980 5448 1992
rect 5500 1980 5506 2032
<< via1 >>
rect 4068 13812 4120 13864
rect 5816 13812 5868 13864
rect 2410 13574 2462 13626
rect 2474 13574 2526 13626
rect 2538 13574 2590 13626
rect 2602 13574 2654 13626
rect 2666 13574 2718 13626
rect 5331 13574 5383 13626
rect 5395 13574 5447 13626
rect 5459 13574 5511 13626
rect 5523 13574 5575 13626
rect 5587 13574 5639 13626
rect 8252 13574 8304 13626
rect 8316 13574 8368 13626
rect 8380 13574 8432 13626
rect 8444 13574 8496 13626
rect 8508 13574 8560 13626
rect 11173 13574 11225 13626
rect 11237 13574 11289 13626
rect 11301 13574 11353 13626
rect 11365 13574 11417 13626
rect 11429 13574 11481 13626
rect 6552 13404 6604 13456
rect 4896 13311 4948 13320
rect 4896 13277 4905 13311
rect 4905 13277 4939 13311
rect 4939 13277 4948 13311
rect 4896 13268 4948 13277
rect 5632 13311 5684 13320
rect 5632 13277 5641 13311
rect 5641 13277 5675 13311
rect 5675 13277 5684 13311
rect 5632 13268 5684 13277
rect 7288 13336 7340 13388
rect 6460 13311 6512 13320
rect 6460 13277 6469 13311
rect 6469 13277 6503 13311
rect 6503 13277 6512 13311
rect 6460 13268 6512 13277
rect 6736 13311 6788 13320
rect 6736 13277 6745 13311
rect 6745 13277 6779 13311
rect 6779 13277 6788 13311
rect 6736 13268 6788 13277
rect 13544 13336 13596 13388
rect 5908 13132 5960 13184
rect 12256 13175 12308 13184
rect 12256 13141 12265 13175
rect 12265 13141 12299 13175
rect 12299 13141 12308 13175
rect 12256 13132 12308 13141
rect 3070 13030 3122 13082
rect 3134 13030 3186 13082
rect 3198 13030 3250 13082
rect 3262 13030 3314 13082
rect 3326 13030 3378 13082
rect 5991 13030 6043 13082
rect 6055 13030 6107 13082
rect 6119 13030 6171 13082
rect 6183 13030 6235 13082
rect 6247 13030 6299 13082
rect 8912 13030 8964 13082
rect 8976 13030 9028 13082
rect 9040 13030 9092 13082
rect 9104 13030 9156 13082
rect 9168 13030 9220 13082
rect 11833 13030 11885 13082
rect 11897 13030 11949 13082
rect 11961 13030 12013 13082
rect 12025 13030 12077 13082
rect 12089 13030 12141 13082
rect 5908 12928 5960 12980
rect 4896 12903 4948 12912
rect 4896 12869 4930 12903
rect 4930 12869 4948 12903
rect 4896 12860 4948 12869
rect 6736 12835 6788 12844
rect 6736 12801 6770 12835
rect 6770 12801 6788 12835
rect 6736 12792 6788 12801
rect 7932 12835 7984 12844
rect 7932 12801 7941 12835
rect 7941 12801 7975 12835
rect 7975 12801 7984 12835
rect 7932 12792 7984 12801
rect 4620 12767 4672 12776
rect 4620 12733 4629 12767
rect 4629 12733 4663 12767
rect 4663 12733 4672 12767
rect 4620 12724 4672 12733
rect 6460 12767 6512 12776
rect 6460 12733 6469 12767
rect 6469 12733 6503 12767
rect 6503 12733 6512 12767
rect 6460 12724 6512 12733
rect 4528 12631 4580 12640
rect 4528 12597 4537 12631
rect 4537 12597 4571 12631
rect 4571 12597 4580 12631
rect 4528 12588 4580 12597
rect 8116 12631 8168 12640
rect 8116 12597 8125 12631
rect 8125 12597 8159 12631
rect 8159 12597 8168 12631
rect 8116 12588 8168 12597
rect 2410 12486 2462 12538
rect 2474 12486 2526 12538
rect 2538 12486 2590 12538
rect 2602 12486 2654 12538
rect 2666 12486 2718 12538
rect 5331 12486 5383 12538
rect 5395 12486 5447 12538
rect 5459 12486 5511 12538
rect 5523 12486 5575 12538
rect 5587 12486 5639 12538
rect 8252 12486 8304 12538
rect 8316 12486 8368 12538
rect 8380 12486 8432 12538
rect 8444 12486 8496 12538
rect 8508 12486 8560 12538
rect 11173 12486 11225 12538
rect 11237 12486 11289 12538
rect 11301 12486 11353 12538
rect 11365 12486 11417 12538
rect 11429 12486 11481 12538
rect 4620 12384 4672 12436
rect 5724 12427 5776 12436
rect 5724 12393 5733 12427
rect 5733 12393 5767 12427
rect 5767 12393 5776 12427
rect 5724 12384 5776 12393
rect 7932 12384 7984 12436
rect 8024 12291 8076 12300
rect 8024 12257 8033 12291
rect 8033 12257 8067 12291
rect 8067 12257 8076 12291
rect 8024 12248 8076 12257
rect 4436 12180 4488 12232
rect 6460 12180 6512 12232
rect 6828 12180 6880 12232
rect 7288 12223 7340 12232
rect 7288 12189 7297 12223
rect 7297 12189 7331 12223
rect 7331 12189 7340 12223
rect 7288 12180 7340 12189
rect 7656 12223 7708 12232
rect 7656 12189 7665 12223
rect 7665 12189 7699 12223
rect 7699 12189 7708 12223
rect 7656 12180 7708 12189
rect 8116 12223 8168 12232
rect 8116 12189 8125 12223
rect 8125 12189 8159 12223
rect 8159 12189 8168 12223
rect 8116 12180 8168 12189
rect 8668 12223 8720 12232
rect 8668 12189 8677 12223
rect 8677 12189 8711 12223
rect 8711 12189 8720 12223
rect 8668 12180 8720 12189
rect 6368 12112 6420 12164
rect 3070 11942 3122 11994
rect 3134 11942 3186 11994
rect 3198 11942 3250 11994
rect 3262 11942 3314 11994
rect 3326 11942 3378 11994
rect 5991 11942 6043 11994
rect 6055 11942 6107 11994
rect 6119 11942 6171 11994
rect 6183 11942 6235 11994
rect 6247 11942 6299 11994
rect 8912 11942 8964 11994
rect 8976 11942 9028 11994
rect 9040 11942 9092 11994
rect 9104 11942 9156 11994
rect 9168 11942 9220 11994
rect 11833 11942 11885 11994
rect 11897 11942 11949 11994
rect 11961 11942 12013 11994
rect 12025 11942 12077 11994
rect 12089 11942 12141 11994
rect 7656 11840 7708 11892
rect 4620 11704 4672 11756
rect 6368 11747 6420 11756
rect 6368 11713 6377 11747
rect 6377 11713 6411 11747
rect 6411 11713 6420 11747
rect 6368 11704 6420 11713
rect 8668 11840 8720 11892
rect 8852 11747 8904 11756
rect 8852 11713 8861 11747
rect 8861 11713 8895 11747
rect 8895 11713 8904 11747
rect 8852 11704 8904 11713
rect 6828 11636 6880 11688
rect 6920 11500 6972 11552
rect 2410 11398 2462 11450
rect 2474 11398 2526 11450
rect 2538 11398 2590 11450
rect 2602 11398 2654 11450
rect 2666 11398 2718 11450
rect 5331 11398 5383 11450
rect 5395 11398 5447 11450
rect 5459 11398 5511 11450
rect 5523 11398 5575 11450
rect 5587 11398 5639 11450
rect 8252 11398 8304 11450
rect 8316 11398 8368 11450
rect 8380 11398 8432 11450
rect 8444 11398 8496 11450
rect 8508 11398 8560 11450
rect 11173 11398 11225 11450
rect 11237 11398 11289 11450
rect 11301 11398 11353 11450
rect 11365 11398 11417 11450
rect 11429 11398 11481 11450
rect 6368 11339 6420 11348
rect 6368 11305 6377 11339
rect 6377 11305 6411 11339
rect 6411 11305 6420 11339
rect 6368 11296 6420 11305
rect 6920 11296 6972 11348
rect 8852 11296 8904 11348
rect 4620 11160 4672 11212
rect 6552 11160 6604 11212
rect 6368 11092 6420 11144
rect 6828 11092 6880 11144
rect 3070 10854 3122 10906
rect 3134 10854 3186 10906
rect 3198 10854 3250 10906
rect 3262 10854 3314 10906
rect 3326 10854 3378 10906
rect 5991 10854 6043 10906
rect 6055 10854 6107 10906
rect 6119 10854 6171 10906
rect 6183 10854 6235 10906
rect 6247 10854 6299 10906
rect 8912 10854 8964 10906
rect 8976 10854 9028 10906
rect 9040 10854 9092 10906
rect 9104 10854 9156 10906
rect 9168 10854 9220 10906
rect 11833 10854 11885 10906
rect 11897 10854 11949 10906
rect 11961 10854 12013 10906
rect 12025 10854 12077 10906
rect 12089 10854 12141 10906
rect 4620 10752 4672 10804
rect 4068 10659 4120 10668
rect 4068 10625 4102 10659
rect 4102 10625 4120 10659
rect 4068 10616 4120 10625
rect 3608 10412 3660 10464
rect 5172 10455 5224 10464
rect 5172 10421 5181 10455
rect 5181 10421 5215 10455
rect 5215 10421 5224 10455
rect 5172 10412 5224 10421
rect 5724 10455 5776 10464
rect 5724 10421 5733 10455
rect 5733 10421 5767 10455
rect 5767 10421 5776 10455
rect 5724 10412 5776 10421
rect 2410 10310 2462 10362
rect 2474 10310 2526 10362
rect 2538 10310 2590 10362
rect 2602 10310 2654 10362
rect 2666 10310 2718 10362
rect 5331 10310 5383 10362
rect 5395 10310 5447 10362
rect 5459 10310 5511 10362
rect 5523 10310 5575 10362
rect 5587 10310 5639 10362
rect 8252 10310 8304 10362
rect 8316 10310 8368 10362
rect 8380 10310 8432 10362
rect 8444 10310 8496 10362
rect 8508 10310 8560 10362
rect 11173 10310 11225 10362
rect 11237 10310 11289 10362
rect 11301 10310 11353 10362
rect 11365 10310 11417 10362
rect 11429 10310 11481 10362
rect 4068 10251 4120 10260
rect 4068 10217 4077 10251
rect 4077 10217 4111 10251
rect 4111 10217 4120 10251
rect 4068 10208 4120 10217
rect 5172 10208 5224 10260
rect 1400 10004 1452 10056
rect 4712 10047 4764 10056
rect 4712 10013 4721 10047
rect 4721 10013 4755 10047
rect 4755 10013 4764 10047
rect 4712 10004 4764 10013
rect 5080 10047 5132 10056
rect 5080 10013 5089 10047
rect 5089 10013 5123 10047
rect 5123 10013 5132 10047
rect 5080 10004 5132 10013
rect 6368 10004 6420 10056
rect 2780 9936 2832 9988
rect 5908 9936 5960 9988
rect 6920 9979 6972 9988
rect 6920 9945 6954 9979
rect 6954 9945 6972 9979
rect 6920 9936 6972 9945
rect 4804 9911 4856 9920
rect 4804 9877 4813 9911
rect 4813 9877 4847 9911
rect 4847 9877 4856 9911
rect 4804 9868 4856 9877
rect 7380 9868 7432 9920
rect 8024 9911 8076 9920
rect 8024 9877 8033 9911
rect 8033 9877 8067 9911
rect 8067 9877 8076 9911
rect 8024 9868 8076 9877
rect 3070 9766 3122 9818
rect 3134 9766 3186 9818
rect 3198 9766 3250 9818
rect 3262 9766 3314 9818
rect 3326 9766 3378 9818
rect 5991 9766 6043 9818
rect 6055 9766 6107 9818
rect 6119 9766 6171 9818
rect 6183 9766 6235 9818
rect 6247 9766 6299 9818
rect 8912 9766 8964 9818
rect 8976 9766 9028 9818
rect 9040 9766 9092 9818
rect 9104 9766 9156 9818
rect 9168 9766 9220 9818
rect 11833 9766 11885 9818
rect 11897 9766 11949 9818
rect 11961 9766 12013 9818
rect 12025 9766 12077 9818
rect 12089 9766 12141 9818
rect 4712 9707 4764 9716
rect 4712 9673 4721 9707
rect 4721 9673 4755 9707
rect 4755 9673 4764 9707
rect 4712 9664 4764 9673
rect 8024 9664 8076 9716
rect 1400 9528 1452 9580
rect 3792 9596 3844 9648
rect 5080 9639 5132 9648
rect 5080 9605 5114 9639
rect 5114 9605 5132 9639
rect 5080 9596 5132 9605
rect 3608 9571 3660 9580
rect 3608 9537 3642 9571
rect 3642 9537 3660 9571
rect 3608 9528 3660 9537
rect 4620 9528 4672 9580
rect 5908 9528 5960 9580
rect 6920 9571 6972 9580
rect 6920 9537 6929 9571
rect 6929 9537 6963 9571
rect 6963 9537 6972 9571
rect 6920 9528 6972 9537
rect 7380 9571 7432 9580
rect 7380 9537 7389 9571
rect 7389 9537 7423 9571
rect 7423 9537 7432 9571
rect 7380 9528 7432 9537
rect 2780 9503 2832 9512
rect 2780 9469 2789 9503
rect 2789 9469 2823 9503
rect 2823 9469 2832 9503
rect 2780 9460 2832 9469
rect 7196 9503 7248 9512
rect 7196 9469 7205 9503
rect 7205 9469 7239 9503
rect 7239 9469 7248 9503
rect 7196 9460 7248 9469
rect 5908 9324 5960 9376
rect 7472 9367 7524 9376
rect 7472 9333 7481 9367
rect 7481 9333 7515 9367
rect 7515 9333 7524 9367
rect 7472 9324 7524 9333
rect 2410 9222 2462 9274
rect 2474 9222 2526 9274
rect 2538 9222 2590 9274
rect 2602 9222 2654 9274
rect 2666 9222 2718 9274
rect 5331 9222 5383 9274
rect 5395 9222 5447 9274
rect 5459 9222 5511 9274
rect 5523 9222 5575 9274
rect 5587 9222 5639 9274
rect 8252 9222 8304 9274
rect 8316 9222 8368 9274
rect 8380 9222 8432 9274
rect 8444 9222 8496 9274
rect 8508 9222 8560 9274
rect 11173 9222 11225 9274
rect 11237 9222 11289 9274
rect 11301 9222 11353 9274
rect 11365 9222 11417 9274
rect 11429 9222 11481 9274
rect 7196 9120 7248 9172
rect 7472 9120 7524 9172
rect 3792 9027 3844 9036
rect 3792 8993 3801 9027
rect 3801 8993 3835 9027
rect 3835 8993 3844 9027
rect 3792 8984 3844 8993
rect 1860 8959 1912 8968
rect 1860 8925 1869 8959
rect 1869 8925 1903 8959
rect 1903 8925 1912 8959
rect 1860 8916 1912 8925
rect 2136 8959 2188 8968
rect 2136 8925 2145 8959
rect 2145 8925 2179 8959
rect 2179 8925 2188 8959
rect 2136 8916 2188 8925
rect 6920 8959 6972 8968
rect 6920 8925 6929 8959
rect 6929 8925 6963 8959
rect 6963 8925 6972 8959
rect 6920 8916 6972 8925
rect 7196 8959 7248 8968
rect 7196 8925 7205 8959
rect 7205 8925 7239 8959
rect 7239 8925 7248 8959
rect 7196 8916 7248 8925
rect 7932 8959 7984 8968
rect 7932 8925 7941 8959
rect 7941 8925 7975 8959
rect 7975 8925 7984 8959
rect 7932 8916 7984 8925
rect 3884 8848 3936 8900
rect 5356 8848 5408 8900
rect 5724 8891 5776 8900
rect 5724 8857 5758 8891
rect 5758 8857 5776 8891
rect 5724 8848 5776 8857
rect 6368 8848 6420 8900
rect 7748 8891 7800 8900
rect 7748 8857 7757 8891
rect 7757 8857 7791 8891
rect 7791 8857 7800 8891
rect 7748 8848 7800 8857
rect 8760 8916 8812 8968
rect 9312 8916 9364 8968
rect 9956 8848 10008 8900
rect 3792 8780 3844 8832
rect 5172 8823 5224 8832
rect 5172 8789 5181 8823
rect 5181 8789 5215 8823
rect 5215 8789 5224 8823
rect 5172 8780 5224 8789
rect 3070 8678 3122 8730
rect 3134 8678 3186 8730
rect 3198 8678 3250 8730
rect 3262 8678 3314 8730
rect 3326 8678 3378 8730
rect 5991 8678 6043 8730
rect 6055 8678 6107 8730
rect 6119 8678 6171 8730
rect 6183 8678 6235 8730
rect 6247 8678 6299 8730
rect 8912 8678 8964 8730
rect 8976 8678 9028 8730
rect 9040 8678 9092 8730
rect 9104 8678 9156 8730
rect 9168 8678 9220 8730
rect 11833 8678 11885 8730
rect 11897 8678 11949 8730
rect 11961 8678 12013 8730
rect 12025 8678 12077 8730
rect 12089 8678 12141 8730
rect 3976 8576 4028 8628
rect 1860 8551 1912 8560
rect 1860 8517 1894 8551
rect 1894 8517 1912 8551
rect 1860 8508 1912 8517
rect 4160 8508 4212 8560
rect 3332 8483 3384 8492
rect 3332 8449 3341 8483
rect 3341 8449 3375 8483
rect 3375 8449 3384 8483
rect 3332 8440 3384 8449
rect 1400 8372 1452 8424
rect 3792 8483 3844 8492
rect 3792 8449 3801 8483
rect 3801 8449 3835 8483
rect 3835 8449 3844 8483
rect 3792 8440 3844 8449
rect 3884 8483 3936 8492
rect 3884 8449 3893 8483
rect 3893 8449 3927 8483
rect 3927 8449 3936 8483
rect 3884 8440 3936 8449
rect 3976 8483 4028 8492
rect 3976 8449 3985 8483
rect 3985 8449 4019 8483
rect 4019 8449 4028 8483
rect 3976 8440 4028 8449
rect 4804 8576 4856 8628
rect 5172 8576 5224 8628
rect 5356 8576 5408 8628
rect 5908 8576 5960 8628
rect 4068 8279 4120 8288
rect 4068 8245 4077 8279
rect 4077 8245 4111 8279
rect 4111 8245 4120 8279
rect 4068 8236 4120 8245
rect 4528 8236 4580 8288
rect 4896 8483 4948 8492
rect 4896 8449 4905 8483
rect 4905 8449 4939 8483
rect 4939 8449 4948 8483
rect 4896 8440 4948 8449
rect 5724 8551 5776 8560
rect 5724 8517 5733 8551
rect 5733 8517 5767 8551
rect 5767 8517 5776 8551
rect 5724 8508 5776 8517
rect 6920 8576 6972 8628
rect 7932 8619 7984 8628
rect 7932 8585 7941 8619
rect 7941 8585 7975 8619
rect 7975 8585 7984 8619
rect 7932 8576 7984 8585
rect 8760 8576 8812 8628
rect 9956 8619 10008 8628
rect 9956 8585 9965 8619
rect 9965 8585 9999 8619
rect 9999 8585 10008 8619
rect 9956 8576 10008 8585
rect 7840 8483 7892 8492
rect 7840 8449 7849 8483
rect 7849 8449 7883 8483
rect 7883 8449 7892 8483
rect 7840 8440 7892 8449
rect 4712 8347 4764 8356
rect 4712 8313 4721 8347
rect 4721 8313 4755 8347
rect 4755 8313 4764 8347
rect 4712 8304 4764 8313
rect 4988 8304 5040 8356
rect 10048 8483 10100 8492
rect 10048 8449 10057 8483
rect 10057 8449 10091 8483
rect 10091 8449 10100 8483
rect 10048 8440 10100 8449
rect 5908 8279 5960 8288
rect 5908 8245 5917 8279
rect 5917 8245 5951 8279
rect 5951 8245 5960 8279
rect 5908 8236 5960 8245
rect 6276 8236 6328 8288
rect 6368 8236 6420 8288
rect 8576 8236 8628 8288
rect 2410 8134 2462 8186
rect 2474 8134 2526 8186
rect 2538 8134 2590 8186
rect 2602 8134 2654 8186
rect 2666 8134 2718 8186
rect 5331 8134 5383 8186
rect 5395 8134 5447 8186
rect 5459 8134 5511 8186
rect 5523 8134 5575 8186
rect 5587 8134 5639 8186
rect 8252 8134 8304 8186
rect 8316 8134 8368 8186
rect 8380 8134 8432 8186
rect 8444 8134 8496 8186
rect 8508 8134 8560 8186
rect 11173 8134 11225 8186
rect 11237 8134 11289 8186
rect 11301 8134 11353 8186
rect 11365 8134 11417 8186
rect 11429 8134 11481 8186
rect 3332 8032 3384 8084
rect 3976 8032 4028 8084
rect 4896 8032 4948 8084
rect 10048 8032 10100 8084
rect 1400 7939 1452 7948
rect 1400 7905 1409 7939
rect 1409 7905 1443 7939
rect 1443 7905 1452 7939
rect 1400 7896 1452 7905
rect 7104 7896 7156 7948
rect 8576 7896 8628 7948
rect 2136 7828 2188 7880
rect 3884 7871 3936 7880
rect 3884 7837 3893 7871
rect 3893 7837 3927 7871
rect 3927 7837 3936 7871
rect 3884 7828 3936 7837
rect 4068 7871 4120 7880
rect 4068 7837 4077 7871
rect 4077 7837 4111 7871
rect 4111 7837 4120 7871
rect 4068 7828 4120 7837
rect 4528 7871 4580 7880
rect 4528 7837 4537 7871
rect 4537 7837 4571 7871
rect 4571 7837 4580 7871
rect 4528 7828 4580 7837
rect 5816 7871 5868 7880
rect 5816 7837 5825 7871
rect 5825 7837 5859 7871
rect 5859 7837 5868 7871
rect 5816 7828 5868 7837
rect 7748 7828 7800 7880
rect 8116 7871 8168 7880
rect 8116 7837 8125 7871
rect 8125 7837 8159 7871
rect 8159 7837 8168 7871
rect 8116 7828 8168 7837
rect 4620 7760 4672 7812
rect 4804 7760 4856 7812
rect 6276 7760 6328 7812
rect 7656 7803 7708 7812
rect 7656 7769 7665 7803
rect 7665 7769 7699 7803
rect 7699 7769 7708 7803
rect 7656 7760 7708 7769
rect 9312 7760 9364 7812
rect 4344 7692 4396 7744
rect 5080 7735 5132 7744
rect 5080 7701 5089 7735
rect 5089 7701 5123 7735
rect 5123 7701 5132 7735
rect 5080 7692 5132 7701
rect 5356 7692 5408 7744
rect 3070 7590 3122 7642
rect 3134 7590 3186 7642
rect 3198 7590 3250 7642
rect 3262 7590 3314 7642
rect 3326 7590 3378 7642
rect 5991 7590 6043 7642
rect 6055 7590 6107 7642
rect 6119 7590 6171 7642
rect 6183 7590 6235 7642
rect 6247 7590 6299 7642
rect 8912 7590 8964 7642
rect 8976 7590 9028 7642
rect 9040 7590 9092 7642
rect 9104 7590 9156 7642
rect 9168 7590 9220 7642
rect 11833 7590 11885 7642
rect 11897 7590 11949 7642
rect 11961 7590 12013 7642
rect 12025 7590 12077 7642
rect 12089 7590 12141 7642
rect 1400 7488 1452 7540
rect 4804 7488 4856 7540
rect 5908 7488 5960 7540
rect 7840 7488 7892 7540
rect 5172 7420 5224 7472
rect 5356 7420 5408 7472
rect 4528 7352 4580 7404
rect 4988 7352 5040 7404
rect 7196 7420 7248 7472
rect 4436 7327 4488 7336
rect 4436 7293 4445 7327
rect 4445 7293 4479 7327
rect 4479 7293 4488 7327
rect 4436 7284 4488 7293
rect 6368 7395 6420 7404
rect 6368 7361 6377 7395
rect 6377 7361 6411 7395
rect 6411 7361 6420 7395
rect 6368 7352 6420 7361
rect 7748 7352 7800 7404
rect 8024 7352 8076 7404
rect 8852 7352 8904 7404
rect 9588 7352 9640 7404
rect 11060 7352 11112 7404
rect 8576 7284 8628 7336
rect 8668 7327 8720 7336
rect 8668 7293 8677 7327
rect 8677 7293 8711 7327
rect 8711 7293 8720 7327
rect 8668 7284 8720 7293
rect 8760 7327 8812 7336
rect 8760 7293 8769 7327
rect 8769 7293 8803 7327
rect 8803 7293 8812 7327
rect 8760 7284 8812 7293
rect 2228 7191 2280 7200
rect 2228 7157 2237 7191
rect 2237 7157 2271 7191
rect 2271 7157 2280 7191
rect 2228 7148 2280 7157
rect 2504 7191 2556 7200
rect 2504 7157 2513 7191
rect 2513 7157 2547 7191
rect 2547 7157 2556 7191
rect 2504 7148 2556 7157
rect 7288 7148 7340 7200
rect 9772 7148 9824 7200
rect 2410 7046 2462 7098
rect 2474 7046 2526 7098
rect 2538 7046 2590 7098
rect 2602 7046 2654 7098
rect 2666 7046 2718 7098
rect 5331 7046 5383 7098
rect 5395 7046 5447 7098
rect 5459 7046 5511 7098
rect 5523 7046 5575 7098
rect 5587 7046 5639 7098
rect 8252 7046 8304 7098
rect 8316 7046 8368 7098
rect 8380 7046 8432 7098
rect 8444 7046 8496 7098
rect 8508 7046 8560 7098
rect 11173 7046 11225 7098
rect 11237 7046 11289 7098
rect 11301 7046 11353 7098
rect 11365 7046 11417 7098
rect 11429 7046 11481 7098
rect 4068 6944 4120 6996
rect 6368 6944 6420 6996
rect 8668 6944 8720 6996
rect 3700 6876 3752 6928
rect 4896 6876 4948 6928
rect 3884 6808 3936 6860
rect 3976 6851 4028 6860
rect 3976 6817 3985 6851
rect 3985 6817 4019 6851
rect 4019 6817 4028 6851
rect 3976 6808 4028 6817
rect 4252 6808 4304 6860
rect 2780 6740 2832 6792
rect 3516 6740 3568 6792
rect 2320 6672 2372 6724
rect 4160 6715 4212 6724
rect 4160 6681 4169 6715
rect 4169 6681 4203 6715
rect 4203 6681 4212 6715
rect 4160 6672 4212 6681
rect 4344 6783 4396 6792
rect 4344 6749 4353 6783
rect 4353 6749 4387 6783
rect 4387 6749 4396 6783
rect 4344 6740 4396 6749
rect 4620 6783 4672 6792
rect 4620 6749 4629 6783
rect 4629 6749 4663 6783
rect 4663 6749 4672 6783
rect 4620 6740 4672 6749
rect 4804 6783 4856 6792
rect 4804 6749 4813 6783
rect 4813 6749 4847 6783
rect 4847 6749 4856 6783
rect 4804 6740 4856 6749
rect 4988 6783 5040 6792
rect 4988 6749 4997 6783
rect 4997 6749 5031 6783
rect 5031 6749 5040 6783
rect 4988 6740 5040 6749
rect 8760 6876 8812 6928
rect 9956 6876 10008 6928
rect 12256 6808 12308 6860
rect 5264 6783 5316 6792
rect 5264 6749 5275 6783
rect 5275 6749 5309 6783
rect 5309 6749 5316 6783
rect 5264 6740 5316 6749
rect 5816 6740 5868 6792
rect 7288 6740 7340 6792
rect 3424 6604 3476 6656
rect 4712 6604 4764 6656
rect 8852 6672 8904 6724
rect 9312 6672 9364 6724
rect 9588 6783 9640 6792
rect 9588 6749 9597 6783
rect 9597 6749 9631 6783
rect 9631 6749 9640 6783
rect 9588 6740 9640 6749
rect 11060 6740 11112 6792
rect 5724 6604 5776 6656
rect 8668 6647 8720 6656
rect 8668 6613 8677 6647
rect 8677 6613 8711 6647
rect 8711 6613 8720 6647
rect 8668 6604 8720 6613
rect 9404 6604 9456 6656
rect 3070 6502 3122 6554
rect 3134 6502 3186 6554
rect 3198 6502 3250 6554
rect 3262 6502 3314 6554
rect 3326 6502 3378 6554
rect 5991 6502 6043 6554
rect 6055 6502 6107 6554
rect 6119 6502 6171 6554
rect 6183 6502 6235 6554
rect 6247 6502 6299 6554
rect 8912 6502 8964 6554
rect 8976 6502 9028 6554
rect 9040 6502 9092 6554
rect 9104 6502 9156 6554
rect 9168 6502 9220 6554
rect 11833 6502 11885 6554
rect 11897 6502 11949 6554
rect 11961 6502 12013 6554
rect 12025 6502 12077 6554
rect 12089 6502 12141 6554
rect 2320 6375 2372 6384
rect 2320 6341 2332 6375
rect 2332 6341 2372 6375
rect 2320 6332 2372 6341
rect 3884 6400 3936 6452
rect 4804 6400 4856 6452
rect 4896 6400 4948 6452
rect 1676 6103 1728 6112
rect 1676 6069 1685 6103
rect 1685 6069 1719 6103
rect 1719 6069 1728 6103
rect 1676 6060 1728 6069
rect 1952 6060 2004 6112
rect 3516 6307 3568 6316
rect 3516 6273 3525 6307
rect 3525 6273 3559 6307
rect 3559 6273 3568 6307
rect 3516 6264 3568 6273
rect 3700 6307 3752 6316
rect 3700 6273 3709 6307
rect 3709 6273 3743 6307
rect 3743 6273 3752 6307
rect 3700 6264 3752 6273
rect 3792 6307 3844 6316
rect 3792 6273 3801 6307
rect 3801 6273 3835 6307
rect 3835 6273 3844 6307
rect 3792 6264 3844 6273
rect 3884 6307 3936 6316
rect 3884 6273 3893 6307
rect 3893 6273 3927 6307
rect 3927 6273 3936 6307
rect 3884 6264 3936 6273
rect 4528 6332 4580 6384
rect 5080 6332 5132 6384
rect 6368 6332 6420 6384
rect 4344 6264 4396 6316
rect 4436 6307 4488 6316
rect 4436 6273 4445 6307
rect 4445 6273 4479 6307
rect 4479 6273 4488 6307
rect 4436 6264 4488 6273
rect 5908 6307 5960 6316
rect 5908 6273 5917 6307
rect 5917 6273 5951 6307
rect 5951 6273 5960 6307
rect 5908 6264 5960 6273
rect 6184 6307 6236 6316
rect 6184 6273 6193 6307
rect 6193 6273 6227 6307
rect 6227 6273 6236 6307
rect 6184 6264 6236 6273
rect 3976 6128 4028 6180
rect 6644 6196 6696 6248
rect 7104 6443 7156 6452
rect 7104 6409 7113 6443
rect 7113 6409 7147 6443
rect 7147 6409 7156 6443
rect 7104 6400 7156 6409
rect 7840 6400 7892 6452
rect 10048 6400 10100 6452
rect 7564 6264 7616 6316
rect 8024 6264 8076 6316
rect 8116 6307 8168 6316
rect 8116 6273 8125 6307
rect 8125 6273 8159 6307
rect 8159 6273 8168 6307
rect 8116 6264 8168 6273
rect 9634 6332 9686 6384
rect 9864 6332 9916 6384
rect 8208 6239 8260 6248
rect 8208 6205 8217 6239
rect 8217 6205 8251 6239
rect 8251 6205 8260 6239
rect 8208 6196 8260 6205
rect 8852 6264 8904 6316
rect 9036 6307 9088 6316
rect 9036 6273 9045 6307
rect 9045 6273 9079 6307
rect 9079 6273 9088 6307
rect 9036 6264 9088 6273
rect 9312 6307 9364 6316
rect 9312 6273 9321 6307
rect 9321 6273 9355 6307
rect 9355 6273 9364 6307
rect 9312 6264 9364 6273
rect 9496 6239 9548 6248
rect 9496 6205 9505 6239
rect 9505 6205 9539 6239
rect 9539 6205 9548 6239
rect 9496 6196 9548 6205
rect 9864 6196 9916 6248
rect 10232 6196 10284 6248
rect 2780 6060 2832 6112
rect 4068 6060 4120 6112
rect 5080 6060 5132 6112
rect 7932 6060 7984 6112
rect 9312 6128 9364 6180
rect 8944 6060 8996 6112
rect 11060 6103 11112 6112
rect 11060 6069 11069 6103
rect 11069 6069 11103 6103
rect 11103 6069 11112 6103
rect 11060 6060 11112 6069
rect 2410 5958 2462 6010
rect 2474 5958 2526 6010
rect 2538 5958 2590 6010
rect 2602 5958 2654 6010
rect 2666 5958 2718 6010
rect 5331 5958 5383 6010
rect 5395 5958 5447 6010
rect 5459 5958 5511 6010
rect 5523 5958 5575 6010
rect 5587 5958 5639 6010
rect 8252 5958 8304 6010
rect 8316 5958 8368 6010
rect 8380 5958 8432 6010
rect 8444 5958 8496 6010
rect 8508 5958 8560 6010
rect 11173 5958 11225 6010
rect 11237 5958 11289 6010
rect 11301 5958 11353 6010
rect 11365 5958 11417 6010
rect 11429 5958 11481 6010
rect 1676 5856 1728 5908
rect 3516 5856 3568 5908
rect 3976 5856 4028 5908
rect 4068 5856 4120 5908
rect 4896 5856 4948 5908
rect 5080 5856 5132 5908
rect 5908 5856 5960 5908
rect 6644 5856 6696 5908
rect 2136 5695 2188 5704
rect 2136 5661 2145 5695
rect 2145 5661 2179 5695
rect 2179 5661 2188 5695
rect 2136 5652 2188 5661
rect 2780 5652 2832 5704
rect 4436 5652 4488 5704
rect 6920 5788 6972 5840
rect 3424 5584 3476 5636
rect 4252 5584 4304 5636
rect 4988 5584 5040 5636
rect 5908 5652 5960 5704
rect 6184 5720 6236 5772
rect 6368 5720 6420 5772
rect 8116 5856 8168 5908
rect 8852 5788 8904 5840
rect 6460 5695 6512 5704
rect 6460 5661 6469 5695
rect 6469 5661 6503 5695
rect 6503 5661 6512 5695
rect 6460 5652 6512 5661
rect 6644 5695 6696 5704
rect 6644 5661 6653 5695
rect 6653 5661 6687 5695
rect 6687 5661 6696 5695
rect 6644 5652 6696 5661
rect 7104 5652 7156 5704
rect 7288 5695 7340 5704
rect 7288 5661 7297 5695
rect 7297 5661 7331 5695
rect 7331 5661 7340 5695
rect 7288 5652 7340 5661
rect 7656 5652 7708 5704
rect 7748 5695 7800 5704
rect 7748 5661 7757 5695
rect 7757 5661 7791 5695
rect 7791 5661 7800 5695
rect 7748 5652 7800 5661
rect 8392 5763 8444 5772
rect 8392 5729 8401 5763
rect 8401 5729 8435 5763
rect 8435 5729 8444 5763
rect 8392 5720 8444 5729
rect 8760 5720 8812 5772
rect 8116 5695 8168 5704
rect 8116 5661 8125 5695
rect 8125 5661 8159 5695
rect 8159 5661 8168 5695
rect 8116 5652 8168 5661
rect 8668 5652 8720 5704
rect 11060 5856 11112 5908
rect 10508 5720 10560 5772
rect 10324 5652 10376 5704
rect 1492 5516 1544 5568
rect 2044 5516 2096 5568
rect 4160 5516 4212 5568
rect 6736 5516 6788 5568
rect 7748 5516 7800 5568
rect 7840 5559 7892 5568
rect 7840 5525 7849 5559
rect 7849 5525 7883 5559
rect 7883 5525 7892 5559
rect 7840 5516 7892 5525
rect 8024 5516 8076 5568
rect 9588 5584 9640 5636
rect 9864 5516 9916 5568
rect 9956 5516 10008 5568
rect 10324 5516 10376 5568
rect 10416 5559 10468 5568
rect 10416 5525 10425 5559
rect 10425 5525 10459 5559
rect 10459 5525 10468 5559
rect 10416 5516 10468 5525
rect 10508 5559 10560 5568
rect 10508 5525 10517 5559
rect 10517 5525 10551 5559
rect 10551 5525 10560 5559
rect 10508 5516 10560 5525
rect 3070 5414 3122 5466
rect 3134 5414 3186 5466
rect 3198 5414 3250 5466
rect 3262 5414 3314 5466
rect 3326 5414 3378 5466
rect 5991 5414 6043 5466
rect 6055 5414 6107 5466
rect 6119 5414 6171 5466
rect 6183 5414 6235 5466
rect 6247 5414 6299 5466
rect 8912 5414 8964 5466
rect 8976 5414 9028 5466
rect 9040 5414 9092 5466
rect 9104 5414 9156 5466
rect 9168 5414 9220 5466
rect 11833 5414 11885 5466
rect 11897 5414 11949 5466
rect 11961 5414 12013 5466
rect 12025 5414 12077 5466
rect 12089 5414 12141 5466
rect 4160 5244 4212 5296
rect 5908 5312 5960 5364
rect 5172 5244 5224 5296
rect 5080 5176 5132 5228
rect 6184 5312 6236 5364
rect 6368 5312 6420 5364
rect 6920 5312 6972 5364
rect 7840 5312 7892 5364
rect 9496 5312 9548 5364
rect 10508 5312 10560 5364
rect 6736 5244 6788 5296
rect 6276 5176 6328 5228
rect 6460 5176 6512 5228
rect 6920 5176 6972 5228
rect 2780 5151 2832 5160
rect 2780 5117 2789 5151
rect 2789 5117 2823 5151
rect 2823 5117 2832 5151
rect 2780 5108 2832 5117
rect 1676 5015 1728 5024
rect 1676 4981 1685 5015
rect 1685 4981 1719 5015
rect 1719 4981 1728 5015
rect 1676 4972 1728 4981
rect 2044 5015 2096 5024
rect 2044 4981 2053 5015
rect 2053 4981 2087 5015
rect 2087 4981 2096 5015
rect 2044 4972 2096 4981
rect 4804 5040 4856 5092
rect 6092 5108 6144 5160
rect 3424 4972 3476 5024
rect 4344 4972 4396 5024
rect 4620 4972 4672 5024
rect 4988 4972 5040 5024
rect 6368 4972 6420 5024
rect 6644 5015 6696 5024
rect 6644 4981 6653 5015
rect 6653 4981 6687 5015
rect 6687 4981 6696 5015
rect 6644 4972 6696 4981
rect 7748 5176 7800 5228
rect 7840 5219 7892 5228
rect 7840 5185 7849 5219
rect 7849 5185 7883 5219
rect 7883 5185 7892 5219
rect 7840 5176 7892 5185
rect 8576 5176 8628 5228
rect 8944 5219 8996 5228
rect 8944 5185 8953 5219
rect 8953 5185 8987 5219
rect 8987 5185 8996 5219
rect 8944 5176 8996 5185
rect 9220 5176 9272 5228
rect 9588 5176 9640 5228
rect 10416 5217 10468 5228
rect 10416 5183 10425 5217
rect 10425 5183 10459 5217
rect 10459 5183 10468 5217
rect 10416 5176 10468 5183
rect 9772 5108 9824 5160
rect 9956 5151 10008 5160
rect 9956 5117 9965 5151
rect 9965 5117 9999 5151
rect 9999 5117 10008 5151
rect 9956 5108 10008 5117
rect 7104 5083 7156 5092
rect 7104 5049 7113 5083
rect 7113 5049 7147 5083
rect 7147 5049 7156 5083
rect 7104 5040 7156 5049
rect 7288 5040 7340 5092
rect 7472 4972 7524 5024
rect 7748 5015 7800 5024
rect 7748 4981 7757 5015
rect 7757 4981 7791 5015
rect 7791 4981 7800 5015
rect 7748 4972 7800 4981
rect 8392 4972 8444 5024
rect 9496 4972 9548 5024
rect 2410 4870 2462 4922
rect 2474 4870 2526 4922
rect 2538 4870 2590 4922
rect 2602 4870 2654 4922
rect 2666 4870 2718 4922
rect 5331 4870 5383 4922
rect 5395 4870 5447 4922
rect 5459 4870 5511 4922
rect 5523 4870 5575 4922
rect 5587 4870 5639 4922
rect 8252 4870 8304 4922
rect 8316 4870 8368 4922
rect 8380 4870 8432 4922
rect 8444 4870 8496 4922
rect 8508 4870 8560 4922
rect 11173 4870 11225 4922
rect 11237 4870 11289 4922
rect 11301 4870 11353 4922
rect 11365 4870 11417 4922
rect 11429 4870 11481 4922
rect 2044 4768 2096 4820
rect 3516 4700 3568 4752
rect 3792 4743 3844 4752
rect 3792 4709 3801 4743
rect 3801 4709 3835 4743
rect 3835 4709 3844 4743
rect 3792 4700 3844 4709
rect 2596 4632 2648 4684
rect 2780 4564 2832 4616
rect 3700 4564 3752 4616
rect 4344 4607 4396 4616
rect 4344 4573 4353 4607
rect 4353 4573 4387 4607
rect 4387 4573 4396 4607
rect 4344 4564 4396 4573
rect 5448 4768 5500 4820
rect 5080 4632 5132 4684
rect 5540 4632 5592 4684
rect 5264 4607 5316 4616
rect 5264 4573 5273 4607
rect 5273 4573 5307 4607
rect 5307 4573 5316 4607
rect 5264 4564 5316 4573
rect 5724 4768 5776 4820
rect 5816 4632 5868 4684
rect 6460 4768 6512 4820
rect 9312 4768 9364 4820
rect 9496 4768 9548 4820
rect 9772 4811 9824 4820
rect 9772 4777 9781 4811
rect 9781 4777 9815 4811
rect 9815 4777 9824 4811
rect 9772 4768 9824 4777
rect 9864 4811 9916 4820
rect 9864 4777 9873 4811
rect 9873 4777 9907 4811
rect 9907 4777 9916 4811
rect 9864 4768 9916 4777
rect 6184 4607 6236 4616
rect 6184 4573 6193 4607
rect 6193 4573 6227 4607
rect 6227 4573 6236 4607
rect 6184 4564 6236 4573
rect 6276 4607 6328 4616
rect 6276 4573 6285 4607
rect 6285 4573 6319 4607
rect 6319 4573 6328 4607
rect 6276 4564 6328 4573
rect 1676 4539 1728 4548
rect 1676 4505 1710 4539
rect 1710 4505 1728 4539
rect 1676 4496 1728 4505
rect 2044 4496 2096 4548
rect 1952 4428 2004 4480
rect 2136 4428 2188 4480
rect 2688 4428 2740 4480
rect 5540 4496 5592 4548
rect 6644 4632 6696 4684
rect 8116 4700 8168 4752
rect 8944 4700 8996 4752
rect 7472 4607 7524 4616
rect 7472 4573 7481 4607
rect 7481 4573 7515 4607
rect 7515 4573 7524 4607
rect 7472 4564 7524 4573
rect 7656 4564 7708 4616
rect 7840 4564 7892 4616
rect 8484 4564 8536 4616
rect 9220 4675 9272 4684
rect 9220 4641 9229 4675
rect 9229 4641 9263 4675
rect 9263 4641 9272 4675
rect 9220 4632 9272 4641
rect 9680 4632 9732 4684
rect 4620 4428 4672 4480
rect 5356 4428 5408 4480
rect 6828 4496 6880 4548
rect 8024 4496 8076 4548
rect 10048 4564 10100 4616
rect 10232 4607 10284 4616
rect 10232 4573 10241 4607
rect 10241 4573 10275 4607
rect 10275 4573 10284 4607
rect 10232 4564 10284 4573
rect 5908 4428 5960 4480
rect 7564 4428 7616 4480
rect 8668 4428 8720 4480
rect 9588 4539 9640 4548
rect 9588 4505 9597 4539
rect 9597 4505 9631 4539
rect 9631 4505 9640 4539
rect 9588 4496 9640 4505
rect 9404 4428 9456 4480
rect 10048 4471 10100 4480
rect 10048 4437 10057 4471
rect 10057 4437 10091 4471
rect 10091 4437 10100 4471
rect 10048 4428 10100 4437
rect 3070 4326 3122 4378
rect 3134 4326 3186 4378
rect 3198 4326 3250 4378
rect 3262 4326 3314 4378
rect 3326 4326 3378 4378
rect 5991 4326 6043 4378
rect 6055 4326 6107 4378
rect 6119 4326 6171 4378
rect 6183 4326 6235 4378
rect 6247 4326 6299 4378
rect 8912 4326 8964 4378
rect 8976 4326 9028 4378
rect 9040 4326 9092 4378
rect 9104 4326 9156 4378
rect 9168 4326 9220 4378
rect 11833 4326 11885 4378
rect 11897 4326 11949 4378
rect 11961 4326 12013 4378
rect 12025 4326 12077 4378
rect 12089 4326 12141 4378
rect 2780 4224 2832 4276
rect 2596 4156 2648 4208
rect 3424 4224 3476 4276
rect 3608 4224 3660 4276
rect 3148 4156 3200 4208
rect 3792 4156 3844 4208
rect 4620 4224 4672 4276
rect 4988 4224 5040 4276
rect 5264 4224 5316 4276
rect 5356 4224 5408 4276
rect 5540 4224 5592 4276
rect 4160 4088 4212 4140
rect 3700 3995 3752 4004
rect 3700 3961 3709 3995
rect 3709 3961 3743 3995
rect 3743 3961 3752 3995
rect 3700 3952 3752 3961
rect 4896 4088 4948 4140
rect 5080 4088 5132 4140
rect 5448 4088 5500 4140
rect 5632 4131 5684 4140
rect 5632 4097 5641 4131
rect 5641 4097 5675 4131
rect 5675 4097 5684 4131
rect 5632 4088 5684 4097
rect 7748 4224 7800 4276
rect 8944 4267 8996 4276
rect 6828 4156 6880 4208
rect 7104 4156 7156 4208
rect 8944 4233 8953 4267
rect 8953 4233 8987 4267
rect 8987 4233 8996 4267
rect 8944 4224 8996 4233
rect 9496 4224 9548 4276
rect 7932 4156 7984 4208
rect 6460 4088 6512 4140
rect 8484 4156 8536 4208
rect 2228 3884 2280 3936
rect 4068 3884 4120 3936
rect 4252 3884 4304 3936
rect 4620 3927 4672 3936
rect 4620 3893 4629 3927
rect 4629 3893 4663 3927
rect 4663 3893 4672 3927
rect 4620 3884 4672 3893
rect 4988 3927 5040 3936
rect 4988 3893 4997 3927
rect 4997 3893 5031 3927
rect 5031 3893 5040 3927
rect 4988 3884 5040 3893
rect 5080 3884 5132 3936
rect 6368 4063 6420 4072
rect 6368 4029 6377 4063
rect 6377 4029 6411 4063
rect 6411 4029 6420 4063
rect 6368 4020 6420 4029
rect 8668 4131 8720 4140
rect 8668 4097 8677 4131
rect 8677 4097 8711 4131
rect 8711 4097 8720 4131
rect 8668 4088 8720 4097
rect 9312 4156 9364 4208
rect 10048 4156 10100 4208
rect 8852 4088 8904 4140
rect 9036 4088 9088 4140
rect 5724 3884 5776 3936
rect 6092 3884 6144 3936
rect 6276 3884 6328 3936
rect 6736 3884 6788 3936
rect 7012 3884 7064 3936
rect 7656 3884 7708 3936
rect 8668 3884 8720 3936
rect 10600 3927 10652 3936
rect 10600 3893 10609 3927
rect 10609 3893 10643 3927
rect 10643 3893 10652 3927
rect 10600 3884 10652 3893
rect 2410 3782 2462 3834
rect 2474 3782 2526 3834
rect 2538 3782 2590 3834
rect 2602 3782 2654 3834
rect 2666 3782 2718 3834
rect 5331 3782 5383 3834
rect 5395 3782 5447 3834
rect 5459 3782 5511 3834
rect 5523 3782 5575 3834
rect 5587 3782 5639 3834
rect 8252 3782 8304 3834
rect 8316 3782 8368 3834
rect 8380 3782 8432 3834
rect 8444 3782 8496 3834
rect 8508 3782 8560 3834
rect 11173 3782 11225 3834
rect 11237 3782 11289 3834
rect 11301 3782 11353 3834
rect 11365 3782 11417 3834
rect 11429 3782 11481 3834
rect 2136 3680 2188 3732
rect 2872 3544 2924 3596
rect 4620 3680 4672 3732
rect 5724 3680 5776 3732
rect 6552 3680 6604 3732
rect 2688 3476 2740 3528
rect 3424 3519 3476 3528
rect 3424 3485 3433 3519
rect 3433 3485 3467 3519
rect 3467 3485 3476 3519
rect 3424 3476 3476 3485
rect 4344 3544 4396 3596
rect 2964 3408 3016 3460
rect 4252 3519 4304 3528
rect 4252 3485 4261 3519
rect 4261 3485 4295 3519
rect 4295 3485 4304 3519
rect 4252 3476 4304 3485
rect 5908 3612 5960 3664
rect 7288 3680 7340 3732
rect 7748 3680 7800 3732
rect 9588 3680 9640 3732
rect 10232 3680 10284 3732
rect 7472 3612 7524 3664
rect 8116 3612 8168 3664
rect 6736 3544 6788 3596
rect 8760 3544 8812 3596
rect 4712 3519 4764 3528
rect 4712 3485 4721 3519
rect 4721 3485 4755 3519
rect 4755 3485 4764 3519
rect 4712 3476 4764 3485
rect 4804 3519 4856 3528
rect 4804 3485 4837 3519
rect 4837 3485 4856 3519
rect 4804 3476 4856 3485
rect 5172 3476 5224 3528
rect 6092 3476 6144 3528
rect 7472 3476 7524 3528
rect 7656 3519 7708 3528
rect 7656 3485 7665 3519
rect 7665 3485 7699 3519
rect 7699 3485 7708 3519
rect 7656 3476 7708 3485
rect 7932 3476 7984 3528
rect 8576 3476 8628 3528
rect 9496 3544 9548 3596
rect 9312 3476 9364 3528
rect 12256 3476 12308 3528
rect 2320 3340 2372 3392
rect 4620 3451 4672 3460
rect 4620 3417 4629 3451
rect 4629 3417 4663 3451
rect 4663 3417 4672 3451
rect 4620 3408 4672 3417
rect 5724 3408 5776 3460
rect 9036 3408 9088 3460
rect 10600 3408 10652 3460
rect 4988 3383 5040 3392
rect 4988 3349 4997 3383
rect 4997 3349 5031 3383
rect 5031 3349 5040 3383
rect 4988 3340 5040 3349
rect 7932 3383 7984 3392
rect 7932 3349 7941 3383
rect 7941 3349 7975 3383
rect 7975 3349 7984 3383
rect 7932 3340 7984 3349
rect 8944 3340 8996 3392
rect 9496 3340 9548 3392
rect 3070 3238 3122 3290
rect 3134 3238 3186 3290
rect 3198 3238 3250 3290
rect 3262 3238 3314 3290
rect 3326 3238 3378 3290
rect 5991 3238 6043 3290
rect 6055 3238 6107 3290
rect 6119 3238 6171 3290
rect 6183 3238 6235 3290
rect 6247 3238 6299 3290
rect 8912 3238 8964 3290
rect 8976 3238 9028 3290
rect 9040 3238 9092 3290
rect 9104 3238 9156 3290
rect 9168 3238 9220 3290
rect 11833 3238 11885 3290
rect 11897 3238 11949 3290
rect 11961 3238 12013 3290
rect 12025 3238 12077 3290
rect 12089 3238 12141 3290
rect 4528 3136 4580 3188
rect 1584 3111 1636 3120
rect 1584 3077 1593 3111
rect 1593 3077 1627 3111
rect 1627 3077 1636 3111
rect 1584 3068 1636 3077
rect 2320 3068 2372 3120
rect 5080 3136 5132 3188
rect 6368 3136 6420 3188
rect 6552 3136 6604 3188
rect 6644 3136 6696 3188
rect 7932 3136 7984 3188
rect 9496 3136 9548 3188
rect 1492 3043 1544 3052
rect 1492 3009 1501 3043
rect 1501 3009 1535 3043
rect 1535 3009 1544 3043
rect 1492 3000 1544 3009
rect 2044 3043 2096 3052
rect 2044 3009 2053 3043
rect 2053 3009 2087 3043
rect 2087 3009 2096 3043
rect 2044 3000 2096 3009
rect 2688 3000 2740 3052
rect 3056 3043 3108 3052
rect 3056 3009 3065 3043
rect 3065 3009 3099 3043
rect 3099 3009 3108 3043
rect 3056 3000 3108 3009
rect 3424 3000 3476 3052
rect 2136 2932 2188 2984
rect 4252 3000 4304 3052
rect 4436 3000 4488 3052
rect 4804 3068 4856 3120
rect 4988 3068 5040 3120
rect 5080 3043 5132 3052
rect 5080 3009 5089 3043
rect 5089 3009 5123 3043
rect 5123 3009 5132 3043
rect 5080 3000 5132 3009
rect 5908 3068 5960 3120
rect 5724 3000 5776 3052
rect 6092 3000 6144 3052
rect 6460 3000 6512 3052
rect 6644 3043 6696 3052
rect 6644 3009 6653 3043
rect 6653 3009 6687 3043
rect 6687 3009 6696 3043
rect 6644 3000 6696 3009
rect 3700 2975 3752 2984
rect 3700 2941 3709 2975
rect 3709 2941 3743 2975
rect 3743 2941 3752 2975
rect 3700 2932 3752 2941
rect 2872 2864 2924 2916
rect 4528 2932 4580 2984
rect 4988 2975 5040 2984
rect 4988 2941 4997 2975
rect 4997 2941 5031 2975
rect 5031 2941 5040 2975
rect 4988 2932 5040 2941
rect 5816 2932 5868 2984
rect 7288 3068 7340 3120
rect 7472 3068 7524 3120
rect 8760 3000 8812 3052
rect 6000 2864 6052 2916
rect 8576 2932 8628 2984
rect 4436 2839 4488 2848
rect 4436 2805 4445 2839
rect 4445 2805 4479 2839
rect 4479 2805 4488 2839
rect 4436 2796 4488 2805
rect 4528 2839 4580 2848
rect 4528 2805 4537 2839
rect 4537 2805 4571 2839
rect 4571 2805 4580 2839
rect 4528 2796 4580 2805
rect 5816 2796 5868 2848
rect 7012 2907 7064 2916
rect 7012 2873 7021 2907
rect 7021 2873 7055 2907
rect 7055 2873 7064 2907
rect 7012 2864 7064 2873
rect 6920 2796 6972 2848
rect 9680 2864 9732 2916
rect 2410 2694 2462 2746
rect 2474 2694 2526 2746
rect 2538 2694 2590 2746
rect 2602 2694 2654 2746
rect 2666 2694 2718 2746
rect 5331 2694 5383 2746
rect 5395 2694 5447 2746
rect 5459 2694 5511 2746
rect 5523 2694 5575 2746
rect 5587 2694 5639 2746
rect 8252 2694 8304 2746
rect 8316 2694 8368 2746
rect 8380 2694 8432 2746
rect 8444 2694 8496 2746
rect 8508 2694 8560 2746
rect 11173 2694 11225 2746
rect 11237 2694 11289 2746
rect 11301 2694 11353 2746
rect 11365 2694 11417 2746
rect 11429 2694 11481 2746
rect 1952 2592 2004 2644
rect 2872 2592 2924 2644
rect 2228 2499 2280 2508
rect 2228 2465 2237 2499
rect 2237 2465 2271 2499
rect 2271 2465 2280 2499
rect 2228 2456 2280 2465
rect 2320 2456 2372 2508
rect 2136 2431 2188 2440
rect 2136 2397 2150 2431
rect 2150 2397 2184 2431
rect 2184 2397 2188 2431
rect 2136 2388 2188 2397
rect 3056 2431 3108 2440
rect 3056 2397 3065 2431
rect 3065 2397 3099 2431
rect 3099 2397 3108 2431
rect 3056 2388 3108 2397
rect 4528 2592 4580 2644
rect 4804 2592 4856 2644
rect 8116 2635 8168 2644
rect 8116 2601 8125 2635
rect 8125 2601 8159 2635
rect 8159 2601 8168 2635
rect 8116 2592 8168 2601
rect 8576 2635 8628 2644
rect 8576 2601 8585 2635
rect 8585 2601 8619 2635
rect 8619 2601 8628 2635
rect 8576 2592 8628 2601
rect 8668 2635 8720 2644
rect 8668 2601 8677 2635
rect 8677 2601 8711 2635
rect 8711 2601 8720 2635
rect 8668 2592 8720 2601
rect 9036 2635 9088 2644
rect 9036 2601 9045 2635
rect 9045 2601 9079 2635
rect 9079 2601 9088 2635
rect 9036 2592 9088 2601
rect 12256 2635 12308 2644
rect 12256 2601 12265 2635
rect 12265 2601 12299 2635
rect 12299 2601 12308 2635
rect 12256 2592 12308 2601
rect 5448 2524 5500 2576
rect 6092 2524 6144 2576
rect 6736 2499 6788 2508
rect 6736 2465 6745 2499
rect 6745 2465 6779 2499
rect 6779 2465 6788 2499
rect 6736 2456 6788 2465
rect 3884 2388 3936 2440
rect 4160 2388 4212 2440
rect 4436 2388 4488 2440
rect 5724 2388 5776 2440
rect 5816 2431 5868 2440
rect 5816 2397 5825 2431
rect 5825 2397 5859 2431
rect 5859 2397 5868 2431
rect 5816 2388 5868 2397
rect 6000 2388 6052 2440
rect 7012 2431 7064 2440
rect 7012 2397 7035 2431
rect 7035 2397 7064 2431
rect 7012 2388 7064 2397
rect 20 2320 72 2372
rect 4988 2320 5040 2372
rect 3608 2252 3660 2304
rect 3792 2295 3844 2304
rect 3792 2261 3801 2295
rect 3801 2261 3835 2295
rect 3835 2261 3844 2295
rect 3792 2252 3844 2261
rect 4068 2252 4120 2304
rect 5448 2363 5500 2372
rect 5448 2329 5457 2363
rect 5457 2329 5491 2363
rect 5491 2329 5500 2363
rect 5448 2320 5500 2329
rect 9404 2456 9456 2508
rect 9312 2388 9364 2440
rect 9588 2388 9640 2440
rect 9772 2252 9824 2304
rect 12808 2252 12860 2304
rect 3070 2150 3122 2202
rect 3134 2150 3186 2202
rect 3198 2150 3250 2202
rect 3262 2150 3314 2202
rect 3326 2150 3378 2202
rect 5991 2150 6043 2202
rect 6055 2150 6107 2202
rect 6119 2150 6171 2202
rect 6183 2150 6235 2202
rect 6247 2150 6299 2202
rect 8912 2150 8964 2202
rect 8976 2150 9028 2202
rect 9040 2150 9092 2202
rect 9104 2150 9156 2202
rect 9168 2150 9220 2202
rect 11833 2150 11885 2202
rect 11897 2150 11949 2202
rect 11961 2150 12013 2202
rect 12025 2150 12077 2202
rect 12089 2150 12141 2202
rect 3792 2048 3844 2100
rect 5816 2048 5868 2100
rect 4344 1980 4396 2032
rect 5448 1980 5500 2032
<< metal2 >>
rect 13542 15266 13598 16066
rect 4066 15056 4122 15065
rect 4066 14991 4122 15000
rect 4080 13870 4108 14991
rect 4068 13864 4120 13870
rect 4068 13806 4120 13812
rect 5816 13864 5868 13870
rect 5816 13806 5868 13812
rect 2410 13628 2718 13637
rect 2410 13626 2416 13628
rect 2472 13626 2496 13628
rect 2552 13626 2576 13628
rect 2632 13626 2656 13628
rect 2712 13626 2718 13628
rect 2472 13574 2474 13626
rect 2654 13574 2656 13626
rect 2410 13572 2416 13574
rect 2472 13572 2496 13574
rect 2552 13572 2576 13574
rect 2632 13572 2656 13574
rect 2712 13572 2718 13574
rect 2410 13563 2718 13572
rect 5331 13628 5639 13637
rect 5331 13626 5337 13628
rect 5393 13626 5417 13628
rect 5473 13626 5497 13628
rect 5553 13626 5577 13628
rect 5633 13626 5639 13628
rect 5393 13574 5395 13626
rect 5575 13574 5577 13626
rect 5331 13572 5337 13574
rect 5393 13572 5417 13574
rect 5473 13572 5497 13574
rect 5553 13572 5577 13574
rect 5633 13572 5639 13574
rect 5331 13563 5639 13572
rect 4896 13320 4948 13326
rect 4896 13262 4948 13268
rect 5632 13320 5684 13326
rect 5632 13262 5684 13268
rect 3070 13084 3378 13093
rect 3070 13082 3076 13084
rect 3132 13082 3156 13084
rect 3212 13082 3236 13084
rect 3292 13082 3316 13084
rect 3372 13082 3378 13084
rect 3132 13030 3134 13082
rect 3314 13030 3316 13082
rect 3070 13028 3076 13030
rect 3132 13028 3156 13030
rect 3212 13028 3236 13030
rect 3292 13028 3316 13030
rect 3372 13028 3378 13030
rect 3070 13019 3378 13028
rect 4908 12918 4936 13262
rect 4896 12912 4948 12918
rect 4896 12854 4948 12860
rect 5644 12866 5672 13262
rect 5644 12838 5764 12866
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 4528 12640 4580 12646
rect 4528 12582 4580 12588
rect 2410 12540 2718 12549
rect 2410 12538 2416 12540
rect 2472 12538 2496 12540
rect 2552 12538 2576 12540
rect 2632 12538 2656 12540
rect 2712 12538 2718 12540
rect 2472 12486 2474 12538
rect 2654 12486 2656 12538
rect 2410 12484 2416 12486
rect 2472 12484 2496 12486
rect 2552 12484 2576 12486
rect 2632 12484 2656 12486
rect 2712 12484 2718 12486
rect 2410 12475 2718 12484
rect 4540 12434 4568 12582
rect 4632 12442 4660 12718
rect 5331 12540 5639 12549
rect 5331 12538 5337 12540
rect 5393 12538 5417 12540
rect 5473 12538 5497 12540
rect 5553 12538 5577 12540
rect 5633 12538 5639 12540
rect 5393 12486 5395 12538
rect 5575 12486 5577 12538
rect 5331 12484 5337 12486
rect 5393 12484 5417 12486
rect 5473 12484 5497 12486
rect 5553 12484 5577 12486
rect 5633 12484 5639 12486
rect 5331 12475 5639 12484
rect 5736 12442 5764 12838
rect 4448 12406 4568 12434
rect 4620 12436 4672 12442
rect 4448 12238 4476 12406
rect 4620 12378 4672 12384
rect 5724 12436 5776 12442
rect 5724 12378 5776 12384
rect 4436 12232 4488 12238
rect 4436 12174 4488 12180
rect 3070 11996 3378 12005
rect 3070 11994 3076 11996
rect 3132 11994 3156 11996
rect 3212 11994 3236 11996
rect 3292 11994 3316 11996
rect 3372 11994 3378 11996
rect 3132 11942 3134 11994
rect 3314 11942 3316 11994
rect 3070 11940 3076 11942
rect 3132 11940 3156 11942
rect 3212 11940 3236 11942
rect 3292 11940 3316 11942
rect 3372 11940 3378 11942
rect 3070 11931 3378 11940
rect 4632 11762 4660 12378
rect 4620 11756 4672 11762
rect 4620 11698 4672 11704
rect 2410 11452 2718 11461
rect 2410 11450 2416 11452
rect 2472 11450 2496 11452
rect 2552 11450 2576 11452
rect 2632 11450 2656 11452
rect 2712 11450 2718 11452
rect 2472 11398 2474 11450
rect 2654 11398 2656 11450
rect 2410 11396 2416 11398
rect 2472 11396 2496 11398
rect 2552 11396 2576 11398
rect 2632 11396 2656 11398
rect 2712 11396 2718 11398
rect 2410 11387 2718 11396
rect 4632 11218 4660 11698
rect 5331 11452 5639 11461
rect 5331 11450 5337 11452
rect 5393 11450 5417 11452
rect 5473 11450 5497 11452
rect 5553 11450 5577 11452
rect 5633 11450 5639 11452
rect 5393 11398 5395 11450
rect 5575 11398 5577 11450
rect 5331 11396 5337 11398
rect 5393 11396 5417 11398
rect 5473 11396 5497 11398
rect 5553 11396 5577 11398
rect 5633 11396 5639 11398
rect 5331 11387 5639 11396
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 3070 10908 3378 10917
rect 3070 10906 3076 10908
rect 3132 10906 3156 10908
rect 3212 10906 3236 10908
rect 3292 10906 3316 10908
rect 3372 10906 3378 10908
rect 3132 10854 3134 10906
rect 3314 10854 3316 10906
rect 3070 10852 3076 10854
rect 3132 10852 3156 10854
rect 3212 10852 3236 10854
rect 3292 10852 3316 10854
rect 3372 10852 3378 10854
rect 3070 10843 3378 10852
rect 4632 10810 4660 11154
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4068 10668 4120 10674
rect 4068 10610 4120 10616
rect 3608 10464 3660 10470
rect 3608 10406 3660 10412
rect 2410 10364 2718 10373
rect 2410 10362 2416 10364
rect 2472 10362 2496 10364
rect 2552 10362 2576 10364
rect 2632 10362 2656 10364
rect 2712 10362 2718 10364
rect 2472 10310 2474 10362
rect 2654 10310 2656 10362
rect 2410 10308 2416 10310
rect 2472 10308 2496 10310
rect 2552 10308 2576 10310
rect 2632 10308 2656 10310
rect 2712 10308 2718 10310
rect 2410 10299 2718 10308
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1412 9586 1440 9998
rect 2780 9988 2832 9994
rect 2780 9930 2832 9936
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 1412 8430 1440 9522
rect 2792 9518 2820 9930
rect 3070 9820 3378 9829
rect 3070 9818 3076 9820
rect 3132 9818 3156 9820
rect 3212 9818 3236 9820
rect 3292 9818 3316 9820
rect 3372 9818 3378 9820
rect 3132 9766 3134 9818
rect 3314 9766 3316 9818
rect 3070 9764 3076 9766
rect 3132 9764 3156 9766
rect 3212 9764 3236 9766
rect 3292 9764 3316 9766
rect 3372 9764 3378 9766
rect 3070 9755 3378 9764
rect 3620 9586 3648 10406
rect 4080 10266 4108 10610
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 3792 9648 3844 9654
rect 3792 9590 3844 9596
rect 3608 9580 3660 9586
rect 3608 9522 3660 9528
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 2410 9276 2718 9285
rect 2410 9274 2416 9276
rect 2472 9274 2496 9276
rect 2552 9274 2576 9276
rect 2632 9274 2656 9276
rect 2712 9274 2718 9276
rect 2472 9222 2474 9274
rect 2654 9222 2656 9274
rect 2410 9220 2416 9222
rect 2472 9220 2496 9222
rect 2552 9220 2576 9222
rect 2632 9220 2656 9222
rect 2712 9220 2718 9222
rect 2410 9211 2718 9220
rect 3804 9042 3832 9590
rect 4632 9586 4660 10746
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5184 10266 5212 10406
rect 5331 10364 5639 10373
rect 5331 10362 5337 10364
rect 5393 10362 5417 10364
rect 5473 10362 5497 10364
rect 5553 10362 5577 10364
rect 5633 10362 5639 10364
rect 5393 10310 5395 10362
rect 5575 10310 5577 10362
rect 5331 10308 5337 10310
rect 5393 10308 5417 10310
rect 5473 10308 5497 10310
rect 5553 10308 5577 10310
rect 5633 10308 5639 10310
rect 5331 10299 5639 10308
rect 5172 10260 5224 10266
rect 5172 10202 5224 10208
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 4724 9722 4752 9998
rect 4804 9920 4856 9926
rect 4804 9862 4856 9868
rect 4712 9716 4764 9722
rect 4712 9658 4764 9664
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 3792 9036 3844 9042
rect 3792 8978 3844 8984
rect 1860 8968 1912 8974
rect 1860 8910 1912 8916
rect 2136 8968 2188 8974
rect 2136 8910 2188 8916
rect 1872 8566 1900 8910
rect 1860 8560 1912 8566
rect 1860 8502 1912 8508
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1412 7954 1440 8366
rect 1400 7948 1452 7954
rect 1400 7890 1452 7896
rect 1412 7546 1440 7890
rect 2148 7886 2176 8910
rect 3884 8900 3936 8906
rect 3884 8842 3936 8848
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 3070 8732 3378 8741
rect 3070 8730 3076 8732
rect 3132 8730 3156 8732
rect 3212 8730 3236 8732
rect 3292 8730 3316 8732
rect 3372 8730 3378 8732
rect 3132 8678 3134 8730
rect 3314 8678 3316 8730
rect 3070 8676 3076 8678
rect 3132 8676 3156 8678
rect 3212 8676 3236 8678
rect 3292 8676 3316 8678
rect 3372 8676 3378 8678
rect 3070 8667 3378 8676
rect 3804 8498 3832 8774
rect 3896 8498 3924 8842
rect 4816 8634 4844 9862
rect 5092 9654 5120 9998
rect 5080 9648 5132 9654
rect 5080 9590 5132 9596
rect 5331 9276 5639 9285
rect 5331 9274 5337 9276
rect 5393 9274 5417 9276
rect 5473 9274 5497 9276
rect 5553 9274 5577 9276
rect 5633 9274 5639 9276
rect 5393 9222 5395 9274
rect 5575 9222 5577 9274
rect 5331 9220 5337 9222
rect 5393 9220 5417 9222
rect 5473 9220 5497 9222
rect 5553 9220 5577 9222
rect 5633 9220 5639 9222
rect 5331 9211 5639 9220
rect 5736 8906 5764 10406
rect 5356 8900 5408 8906
rect 5356 8842 5408 8848
rect 5724 8900 5776 8906
rect 5724 8842 5776 8848
rect 5172 8832 5224 8838
rect 5172 8774 5224 8780
rect 5184 8634 5212 8774
rect 5368 8634 5396 8842
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 4804 8628 4856 8634
rect 4804 8570 4856 8576
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 3988 8498 4016 8570
rect 4160 8560 4212 8566
rect 4160 8502 4212 8508
rect 5724 8560 5776 8566
rect 5724 8502 5776 8508
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3792 8492 3844 8498
rect 3792 8434 3844 8440
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 3976 8492 4028 8498
rect 3976 8434 4028 8440
rect 2410 8188 2718 8197
rect 2410 8186 2416 8188
rect 2472 8186 2496 8188
rect 2552 8186 2576 8188
rect 2632 8186 2656 8188
rect 2712 8186 2718 8188
rect 2472 8134 2474 8186
rect 2654 8134 2656 8186
rect 2410 8132 2416 8134
rect 2472 8132 2496 8134
rect 2552 8132 2576 8134
rect 2632 8132 2656 8134
rect 2712 8132 2718 8134
rect 2410 8123 2718 8132
rect 3344 8090 3372 8434
rect 3988 8090 4016 8434
rect 4172 8378 4200 8502
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 4172 8350 4476 8378
rect 4068 8288 4120 8294
rect 4120 8236 4292 8242
rect 4068 8230 4292 8236
rect 4080 8214 4292 8230
rect 3332 8084 3384 8090
rect 3332 8026 3384 8032
rect 3976 8084 4028 8090
rect 3976 8026 4028 8032
rect 2136 7880 2188 7886
rect 2136 7822 2188 7828
rect 3884 7880 3936 7886
rect 3884 7822 3936 7828
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 3070 7644 3378 7653
rect 3070 7642 3076 7644
rect 3132 7642 3156 7644
rect 3212 7642 3236 7644
rect 3292 7642 3316 7644
rect 3372 7642 3378 7644
rect 3132 7590 3134 7642
rect 3314 7590 3316 7642
rect 3070 7588 3076 7590
rect 3132 7588 3156 7590
rect 3212 7588 3236 7590
rect 3292 7588 3316 7590
rect 3372 7588 3378 7590
rect 3070 7579 3378 7588
rect 1400 7540 1452 7546
rect 1400 7482 1452 7488
rect 2228 7200 2280 7206
rect 2504 7200 2556 7206
rect 2228 7142 2280 7148
rect 2332 7160 2504 7188
rect 2240 6610 2268 7142
rect 2332 6730 2360 7160
rect 2504 7142 2556 7148
rect 2410 7100 2718 7109
rect 2410 7098 2416 7100
rect 2472 7098 2496 7100
rect 2552 7098 2576 7100
rect 2632 7098 2656 7100
rect 2712 7098 2718 7100
rect 2472 7046 2474 7098
rect 2654 7046 2656 7098
rect 2410 7044 2416 7046
rect 2472 7044 2496 7046
rect 2552 7044 2576 7046
rect 2632 7044 2656 7046
rect 2712 7044 2718 7046
rect 2410 7035 2718 7044
rect 3700 6928 3752 6934
rect 3752 6888 3832 6916
rect 3700 6870 3752 6876
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 3516 6792 3568 6798
rect 3516 6734 3568 6740
rect 2320 6724 2372 6730
rect 2320 6666 2372 6672
rect 2240 6582 2360 6610
rect 2332 6390 2360 6582
rect 2320 6384 2372 6390
rect 2320 6326 2372 6332
rect 2792 6118 2820 6734
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3070 6556 3378 6565
rect 3070 6554 3076 6556
rect 3132 6554 3156 6556
rect 3212 6554 3236 6556
rect 3292 6554 3316 6556
rect 3372 6554 3378 6556
rect 3132 6502 3134 6554
rect 3314 6502 3316 6554
rect 3070 6500 3076 6502
rect 3132 6500 3156 6502
rect 3212 6500 3236 6502
rect 3292 6500 3316 6502
rect 3372 6500 3378 6502
rect 3070 6491 3378 6500
rect 1676 6112 1728 6118
rect 1676 6054 1728 6060
rect 1952 6112 2004 6118
rect 2780 6112 2832 6118
rect 2004 6060 2084 6066
rect 1952 6054 2084 6060
rect 2780 6054 2832 6060
rect 1688 5914 1716 6054
rect 1964 6038 2084 6054
rect 1676 5908 1728 5914
rect 1676 5850 1728 5856
rect 2056 5574 2084 6038
rect 2410 6012 2718 6021
rect 2410 6010 2416 6012
rect 2472 6010 2496 6012
rect 2552 6010 2576 6012
rect 2632 6010 2656 6012
rect 2712 6010 2718 6012
rect 2472 5958 2474 6010
rect 2654 5958 2656 6010
rect 2410 5956 2416 5958
rect 2472 5956 2496 5958
rect 2552 5956 2576 5958
rect 2632 5956 2656 5958
rect 2712 5956 2718 5958
rect 2410 5947 2718 5956
rect 2792 5710 2820 6054
rect 2136 5704 2188 5710
rect 2136 5646 2188 5652
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 1492 5568 1544 5574
rect 1492 5510 1544 5516
rect 2044 5568 2096 5574
rect 2044 5510 2096 5516
rect 1504 4185 1532 5510
rect 1676 5024 1728 5030
rect 1676 4966 1728 4972
rect 2044 5024 2096 5030
rect 2044 4966 2096 4972
rect 1688 4554 1716 4966
rect 2056 4826 2084 4966
rect 2044 4820 2096 4826
rect 2044 4762 2096 4768
rect 1676 4548 1728 4554
rect 1676 4490 1728 4496
rect 2044 4548 2096 4554
rect 2044 4490 2096 4496
rect 1952 4480 2004 4486
rect 1952 4422 2004 4428
rect 1490 4176 1546 4185
rect 1490 4111 1546 4120
rect 1504 3058 1532 4111
rect 1584 3120 1636 3126
rect 1582 3088 1584 3097
rect 1636 3088 1638 3097
rect 1492 3052 1544 3058
rect 1582 3023 1638 3032
rect 1492 2994 1544 3000
rect 1964 2650 1992 4422
rect 2056 3058 2084 4490
rect 2148 4486 2176 5646
rect 2792 5166 2820 5646
rect 3436 5642 3464 6598
rect 3528 6322 3556 6734
rect 3804 6322 3832 6888
rect 3896 6866 3924 7822
rect 4080 7002 4108 7822
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 4264 6866 4292 8214
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 3884 6860 3936 6866
rect 3884 6802 3936 6808
rect 3976 6860 4028 6866
rect 3976 6802 4028 6808
rect 4252 6860 4304 6866
rect 4252 6802 4304 6808
rect 3896 6458 3924 6802
rect 3884 6452 3936 6458
rect 3884 6394 3936 6400
rect 3516 6316 3568 6322
rect 3516 6258 3568 6264
rect 3700 6316 3752 6322
rect 3700 6258 3752 6264
rect 3792 6316 3844 6322
rect 3792 6258 3844 6264
rect 3884 6316 3936 6322
rect 3884 6258 3936 6264
rect 3712 6225 3740 6258
rect 3698 6216 3754 6225
rect 3698 6151 3754 6160
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 3424 5636 3476 5642
rect 3424 5578 3476 5584
rect 3070 5468 3378 5477
rect 3070 5466 3076 5468
rect 3132 5466 3156 5468
rect 3212 5466 3236 5468
rect 3292 5466 3316 5468
rect 3372 5466 3378 5468
rect 3132 5414 3134 5466
rect 3314 5414 3316 5466
rect 3070 5412 3076 5414
rect 3132 5412 3156 5414
rect 3212 5412 3236 5414
rect 3292 5412 3316 5414
rect 3372 5412 3378 5414
rect 3070 5403 3378 5412
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 2410 4924 2718 4933
rect 2410 4922 2416 4924
rect 2472 4922 2496 4924
rect 2552 4922 2576 4924
rect 2632 4922 2656 4924
rect 2712 4922 2718 4924
rect 2472 4870 2474 4922
rect 2654 4870 2656 4922
rect 2410 4868 2416 4870
rect 2472 4868 2496 4870
rect 2552 4868 2576 4870
rect 2632 4868 2656 4870
rect 2712 4868 2718 4870
rect 2410 4859 2718 4868
rect 2596 4684 2648 4690
rect 2596 4626 2648 4632
rect 2136 4480 2188 4486
rect 2136 4422 2188 4428
rect 2608 4214 2636 4626
rect 2792 4622 2820 5102
rect 3424 5024 3476 5030
rect 3424 4966 3476 4972
rect 2780 4616 2832 4622
rect 2780 4558 2832 4564
rect 2688 4480 2740 4486
rect 2688 4422 2740 4428
rect 2596 4208 2648 4214
rect 2596 4150 2648 4156
rect 2228 3936 2280 3942
rect 2700 3924 2728 4422
rect 2792 4298 2820 4558
rect 3070 4380 3378 4389
rect 3070 4378 3076 4380
rect 3132 4378 3156 4380
rect 3212 4378 3236 4380
rect 3292 4378 3316 4380
rect 3372 4378 3378 4380
rect 3132 4326 3134 4378
rect 3314 4326 3316 4378
rect 3070 4324 3076 4326
rect 3132 4324 3156 4326
rect 3212 4324 3236 4326
rect 3292 4324 3316 4326
rect 3372 4324 3378 4326
rect 3070 4315 3378 4324
rect 2792 4282 2912 4298
rect 3436 4282 3464 4966
rect 3528 4758 3556 5850
rect 3896 5137 3924 6258
rect 3988 6186 4016 6802
rect 4160 6724 4212 6730
rect 4160 6666 4212 6672
rect 3976 6180 4028 6186
rect 3976 6122 4028 6128
rect 3988 5914 4016 6122
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 4080 5914 4108 6054
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 4172 5574 4200 6666
rect 4264 5642 4292 6802
rect 4356 6798 4384 7686
rect 4448 7562 4476 8350
rect 4712 8356 4764 8362
rect 4712 8298 4764 8304
rect 4528 8288 4580 8294
rect 4528 8230 4580 8236
rect 4540 7886 4568 8230
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 4620 7812 4672 7818
rect 4620 7754 4672 7760
rect 4448 7534 4568 7562
rect 4540 7410 4568 7534
rect 4528 7404 4580 7410
rect 4528 7346 4580 7352
rect 4436 7336 4488 7342
rect 4436 7278 4488 7284
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 4448 6322 4476 7278
rect 4632 6798 4660 7754
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4724 6662 4752 8298
rect 4908 8090 4936 8434
rect 4988 8356 5040 8362
rect 4988 8298 5040 8304
rect 4896 8084 4948 8090
rect 4896 8026 4948 8032
rect 5000 7970 5028 8298
rect 5331 8188 5639 8197
rect 5331 8186 5337 8188
rect 5393 8186 5417 8188
rect 5473 8186 5497 8188
rect 5553 8186 5577 8188
rect 5633 8186 5639 8188
rect 5393 8134 5395 8186
rect 5575 8134 5577 8186
rect 5331 8132 5337 8134
rect 5393 8132 5417 8134
rect 5473 8132 5497 8134
rect 5553 8132 5577 8134
rect 5633 8132 5639 8134
rect 5331 8123 5639 8132
rect 4908 7942 5028 7970
rect 4804 7812 4856 7818
rect 4804 7754 4856 7760
rect 4816 7546 4844 7754
rect 4804 7540 4856 7546
rect 4804 7482 4856 7488
rect 4908 6934 4936 7942
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 4988 7404 5040 7410
rect 4988 7346 5040 7352
rect 4896 6928 4948 6934
rect 4896 6870 4948 6876
rect 5000 6798 5028 7346
rect 4804 6792 4856 6798
rect 4804 6734 4856 6740
rect 4988 6792 5040 6798
rect 4988 6734 5040 6740
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4816 6458 4844 6734
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 4896 6452 4948 6458
rect 4896 6394 4948 6400
rect 4528 6384 4580 6390
rect 4580 6344 4752 6372
rect 4528 6326 4580 6332
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 4436 6316 4488 6322
rect 4436 6258 4488 6264
rect 4252 5636 4304 5642
rect 4252 5578 4304 5584
rect 4160 5568 4212 5574
rect 4160 5510 4212 5516
rect 4160 5296 4212 5302
rect 4158 5264 4160 5273
rect 4212 5264 4214 5273
rect 4158 5199 4214 5208
rect 3882 5128 3938 5137
rect 3882 5063 3938 5072
rect 3516 4752 3568 4758
rect 3516 4694 3568 4700
rect 3792 4752 3844 4758
rect 3792 4694 3844 4700
rect 3700 4616 3752 4622
rect 3700 4558 3752 4564
rect 2780 4276 2912 4282
rect 2832 4270 2912 4276
rect 2780 4218 2832 4224
rect 2700 3896 2820 3924
rect 2228 3878 2280 3884
rect 2240 3754 2268 3878
rect 2410 3836 2718 3845
rect 2410 3834 2416 3836
rect 2472 3834 2496 3836
rect 2552 3834 2576 3836
rect 2632 3834 2656 3836
rect 2712 3834 2718 3836
rect 2472 3782 2474 3834
rect 2654 3782 2656 3834
rect 2410 3780 2416 3782
rect 2472 3780 2496 3782
rect 2552 3780 2576 3782
rect 2632 3780 2656 3782
rect 2712 3780 2718 3782
rect 2410 3771 2718 3780
rect 2148 3738 2268 3754
rect 2136 3732 2268 3738
rect 2188 3726 2268 3732
rect 2136 3674 2188 3680
rect 2044 3052 2096 3058
rect 2044 2994 2096 3000
rect 2136 2984 2188 2990
rect 2136 2926 2188 2932
rect 1952 2644 2004 2650
rect 1952 2586 2004 2592
rect 2148 2446 2176 2926
rect 2240 2514 2268 3726
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 2320 3392 2372 3398
rect 2320 3334 2372 3340
rect 2332 3126 2360 3334
rect 2320 3120 2372 3126
rect 2320 3062 2372 3068
rect 2332 2514 2360 3062
rect 2700 3058 2728 3470
rect 2792 3448 2820 3896
rect 2884 3602 2912 4270
rect 3424 4276 3476 4282
rect 3424 4218 3476 4224
rect 3608 4276 3660 4282
rect 3608 4218 3660 4224
rect 3148 4208 3200 4214
rect 3054 4176 3110 4185
rect 3110 4156 3148 4162
rect 3110 4150 3200 4156
rect 3110 4134 3188 4150
rect 3054 4111 3110 4120
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 3424 3528 3476 3534
rect 3424 3470 3476 3476
rect 2964 3460 3016 3466
rect 2792 3420 2964 3448
rect 2964 3402 3016 3408
rect 3070 3292 3378 3301
rect 3070 3290 3076 3292
rect 3132 3290 3156 3292
rect 3212 3290 3236 3292
rect 3292 3290 3316 3292
rect 3372 3290 3378 3292
rect 3132 3238 3134 3290
rect 3314 3238 3316 3290
rect 3070 3236 3076 3238
rect 3132 3236 3156 3238
rect 3212 3236 3236 3238
rect 3292 3236 3316 3238
rect 3372 3236 3378 3238
rect 3070 3227 3378 3236
rect 3436 3058 3464 3470
rect 2688 3052 2740 3058
rect 2688 2994 2740 3000
rect 3056 3052 3108 3058
rect 3056 2994 3108 3000
rect 3424 3052 3476 3058
rect 3424 2994 3476 3000
rect 2872 2916 2924 2922
rect 2872 2858 2924 2864
rect 2410 2748 2718 2757
rect 2410 2746 2416 2748
rect 2472 2746 2496 2748
rect 2552 2746 2576 2748
rect 2632 2746 2656 2748
rect 2712 2746 2718 2748
rect 2472 2694 2474 2746
rect 2654 2694 2656 2746
rect 2410 2692 2416 2694
rect 2472 2692 2496 2694
rect 2552 2692 2576 2694
rect 2632 2692 2656 2694
rect 2712 2692 2718 2694
rect 2410 2683 2718 2692
rect 2884 2650 2912 2858
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 2228 2508 2280 2514
rect 2228 2450 2280 2456
rect 2320 2508 2372 2514
rect 2320 2450 2372 2456
rect 3068 2446 3096 2994
rect 2136 2440 2188 2446
rect 2136 2382 2188 2388
rect 3056 2440 3108 2446
rect 3056 2382 3108 2388
rect 20 2372 72 2378
rect 20 2314 72 2320
rect 32 800 60 2314
rect 3620 2310 3648 4218
rect 3712 4010 3740 4558
rect 3804 4214 3832 4694
rect 3792 4208 3844 4214
rect 3792 4150 3844 4156
rect 3700 4004 3752 4010
rect 3700 3946 3752 3952
rect 3700 2984 3752 2990
rect 3752 2944 3832 2972
rect 3700 2926 3752 2932
rect 3804 2310 3832 2944
rect 3896 2446 3924 5063
rect 4172 4146 4200 5199
rect 4356 5030 4384 6258
rect 4448 5710 4476 6258
rect 4436 5704 4488 5710
rect 4436 5646 4488 5652
rect 4344 5024 4396 5030
rect 4344 4966 4396 4972
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 4080 2310 4108 3878
rect 4264 3534 4292 3878
rect 4356 3602 4384 4558
rect 4632 4486 4660 4966
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4632 4282 4660 4422
rect 4620 4276 4672 4282
rect 4620 4218 4672 4224
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4632 3738 4660 3878
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 4344 3596 4396 3602
rect 4344 3538 4396 3544
rect 4252 3528 4304 3534
rect 4252 3470 4304 3476
rect 4264 3058 4292 3470
rect 4252 3052 4304 3058
rect 4252 2994 4304 3000
rect 4158 2816 4214 2825
rect 4158 2751 4214 2760
rect 4172 2446 4200 2751
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 3608 2304 3660 2310
rect 3608 2246 3660 2252
rect 3792 2304 3844 2310
rect 3792 2246 3844 2252
rect 4068 2304 4120 2310
rect 4068 2246 4120 2252
rect 3070 2204 3378 2213
rect 3070 2202 3076 2204
rect 3132 2202 3156 2204
rect 3212 2202 3236 2204
rect 3292 2202 3316 2204
rect 3372 2202 3378 2204
rect 3132 2150 3134 2202
rect 3314 2150 3316 2202
rect 3070 2148 3076 2150
rect 3132 2148 3156 2150
rect 3212 2148 3236 2150
rect 3292 2148 3316 2150
rect 3372 2148 3378 2150
rect 3070 2139 3378 2148
rect 3804 2106 3832 2246
rect 3792 2100 3844 2106
rect 3792 2042 3844 2048
rect 4356 2038 4384 3538
rect 4724 3534 4752 6344
rect 4908 5914 4936 6394
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 5000 5642 5028 6734
rect 5092 6390 5120 7686
rect 5368 7478 5396 7686
rect 5172 7472 5224 7478
rect 5172 7414 5224 7420
rect 5356 7472 5408 7478
rect 5356 7414 5408 7420
rect 5184 6780 5212 7414
rect 5331 7100 5639 7109
rect 5331 7098 5337 7100
rect 5393 7098 5417 7100
rect 5473 7098 5497 7100
rect 5553 7098 5577 7100
rect 5633 7098 5639 7100
rect 5393 7046 5395 7098
rect 5575 7046 5577 7098
rect 5331 7044 5337 7046
rect 5393 7044 5417 7046
rect 5473 7044 5497 7046
rect 5553 7044 5577 7046
rect 5633 7044 5639 7046
rect 5331 7035 5639 7044
rect 5264 6792 5316 6798
rect 5184 6752 5264 6780
rect 5080 6384 5132 6390
rect 5080 6326 5132 6332
rect 5080 6112 5132 6118
rect 5080 6054 5132 6060
rect 5092 5914 5120 6054
rect 5080 5908 5132 5914
rect 5080 5850 5132 5856
rect 4988 5636 5040 5642
rect 4988 5578 5040 5584
rect 5184 5302 5212 6752
rect 5264 6734 5316 6740
rect 5736 6662 5764 8502
rect 5828 7886 5856 13806
rect 8252 13628 8560 13637
rect 8252 13626 8258 13628
rect 8314 13626 8338 13628
rect 8394 13626 8418 13628
rect 8474 13626 8498 13628
rect 8554 13626 8560 13628
rect 8314 13574 8316 13626
rect 8496 13574 8498 13626
rect 8252 13572 8258 13574
rect 8314 13572 8338 13574
rect 8394 13572 8418 13574
rect 8474 13572 8498 13574
rect 8554 13572 8560 13574
rect 8252 13563 8560 13572
rect 11173 13628 11481 13637
rect 11173 13626 11179 13628
rect 11235 13626 11259 13628
rect 11315 13626 11339 13628
rect 11395 13626 11419 13628
rect 11475 13626 11481 13628
rect 11235 13574 11237 13626
rect 11417 13574 11419 13626
rect 11173 13572 11179 13574
rect 11235 13572 11259 13574
rect 11315 13572 11339 13574
rect 11395 13572 11419 13574
rect 11475 13572 11481 13574
rect 11173 13563 11481 13572
rect 6552 13456 6604 13462
rect 6552 13398 6604 13404
rect 6460 13320 6512 13326
rect 6460 13262 6512 13268
rect 5908 13184 5960 13190
rect 5908 13126 5960 13132
rect 5920 12986 5948 13126
rect 5991 13084 6299 13093
rect 5991 13082 5997 13084
rect 6053 13082 6077 13084
rect 6133 13082 6157 13084
rect 6213 13082 6237 13084
rect 6293 13082 6299 13084
rect 6053 13030 6055 13082
rect 6235 13030 6237 13082
rect 5991 13028 5997 13030
rect 6053 13028 6077 13030
rect 6133 13028 6157 13030
rect 6213 13028 6237 13030
rect 6293 13028 6299 13030
rect 5991 13019 6299 13028
rect 5908 12980 5960 12986
rect 5908 12922 5960 12928
rect 6472 12866 6500 13262
rect 6380 12838 6500 12866
rect 6380 12170 6408 12838
rect 6460 12776 6512 12782
rect 6460 12718 6512 12724
rect 6472 12238 6500 12718
rect 6460 12232 6512 12238
rect 6460 12174 6512 12180
rect 6368 12164 6420 12170
rect 6368 12106 6420 12112
rect 5991 11996 6299 12005
rect 5991 11994 5997 11996
rect 6053 11994 6077 11996
rect 6133 11994 6157 11996
rect 6213 11994 6237 11996
rect 6293 11994 6299 11996
rect 6053 11942 6055 11994
rect 6235 11942 6237 11994
rect 5991 11940 5997 11942
rect 6053 11940 6077 11942
rect 6133 11940 6157 11942
rect 6213 11940 6237 11942
rect 6293 11940 6299 11942
rect 5991 11931 6299 11940
rect 6368 11756 6420 11762
rect 6368 11698 6420 11704
rect 6380 11354 6408 11698
rect 6368 11348 6420 11354
rect 6368 11290 6420 11296
rect 6564 11218 6592 13398
rect 13556 13394 13584 15266
rect 7288 13388 7340 13394
rect 7288 13330 7340 13336
rect 13544 13388 13596 13394
rect 13544 13330 13596 13336
rect 6736 13320 6788 13326
rect 6736 13262 6788 13268
rect 6748 12850 6776 13262
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 7300 12238 7328 13330
rect 12256 13184 12308 13190
rect 12256 13126 12308 13132
rect 8912 13084 9220 13093
rect 8912 13082 8918 13084
rect 8974 13082 8998 13084
rect 9054 13082 9078 13084
rect 9134 13082 9158 13084
rect 9214 13082 9220 13084
rect 8974 13030 8976 13082
rect 9156 13030 9158 13082
rect 8912 13028 8918 13030
rect 8974 13028 8998 13030
rect 9054 13028 9078 13030
rect 9134 13028 9158 13030
rect 9214 13028 9220 13030
rect 8912 13019 9220 13028
rect 11833 13084 12141 13093
rect 11833 13082 11839 13084
rect 11895 13082 11919 13084
rect 11975 13082 11999 13084
rect 12055 13082 12079 13084
rect 12135 13082 12141 13084
rect 11895 13030 11897 13082
rect 12077 13030 12079 13082
rect 11833 13028 11839 13030
rect 11895 13028 11919 13030
rect 11975 13028 11999 13030
rect 12055 13028 12079 13030
rect 12135 13028 12141 13030
rect 11833 13019 12141 13028
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 7944 12442 7972 12786
rect 8116 12640 8168 12646
rect 8116 12582 8168 12588
rect 7932 12436 7984 12442
rect 7932 12378 7984 12384
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 7288 12232 7340 12238
rect 7288 12174 7340 12180
rect 7656 12232 7708 12238
rect 7656 12174 7708 12180
rect 6840 11694 6868 12174
rect 7668 11898 7696 12174
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 6552 11212 6604 11218
rect 6552 11154 6604 11160
rect 6840 11150 6868 11630
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 6932 11354 6960 11494
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 6368 11144 6420 11150
rect 6368 11086 6420 11092
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 5991 10908 6299 10917
rect 5991 10906 5997 10908
rect 6053 10906 6077 10908
rect 6133 10906 6157 10908
rect 6213 10906 6237 10908
rect 6293 10906 6299 10908
rect 6053 10854 6055 10906
rect 6235 10854 6237 10906
rect 5991 10852 5997 10854
rect 6053 10852 6077 10854
rect 6133 10852 6157 10854
rect 6213 10852 6237 10854
rect 6293 10852 6299 10854
rect 5991 10843 6299 10852
rect 6380 10062 6408 11086
rect 6368 10056 6420 10062
rect 6368 9998 6420 10004
rect 8036 10010 8064 12242
rect 8128 12238 8156 12582
rect 8252 12540 8560 12549
rect 8252 12538 8258 12540
rect 8314 12538 8338 12540
rect 8394 12538 8418 12540
rect 8474 12538 8498 12540
rect 8554 12538 8560 12540
rect 8314 12486 8316 12538
rect 8496 12486 8498 12538
rect 8252 12484 8258 12486
rect 8314 12484 8338 12486
rect 8394 12484 8418 12486
rect 8474 12484 8498 12486
rect 8554 12484 8560 12486
rect 8252 12475 8560 12484
rect 11173 12540 11481 12549
rect 11173 12538 11179 12540
rect 11235 12538 11259 12540
rect 11315 12538 11339 12540
rect 11395 12538 11419 12540
rect 11475 12538 11481 12540
rect 11235 12486 11237 12538
rect 11417 12486 11419 12538
rect 11173 12484 11179 12486
rect 11235 12484 11259 12486
rect 11315 12484 11339 12486
rect 11395 12484 11419 12486
rect 11475 12484 11481 12486
rect 11173 12475 11481 12484
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 8680 11898 8708 12174
rect 8912 11996 9220 12005
rect 8912 11994 8918 11996
rect 8974 11994 8998 11996
rect 9054 11994 9078 11996
rect 9134 11994 9158 11996
rect 9214 11994 9220 11996
rect 8974 11942 8976 11994
rect 9156 11942 9158 11994
rect 8912 11940 8918 11942
rect 8974 11940 8998 11942
rect 9054 11940 9078 11942
rect 9134 11940 9158 11942
rect 9214 11940 9220 11942
rect 8912 11931 9220 11940
rect 11833 11996 12141 12005
rect 11833 11994 11839 11996
rect 11895 11994 11919 11996
rect 11975 11994 11999 11996
rect 12055 11994 12079 11996
rect 12135 11994 12141 11996
rect 11895 11942 11897 11994
rect 12077 11942 12079 11994
rect 11833 11940 11839 11942
rect 11895 11940 11919 11942
rect 11975 11940 11999 11942
rect 12055 11940 12079 11942
rect 12135 11940 12141 11942
rect 11833 11931 12141 11940
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 8252 11452 8560 11461
rect 8252 11450 8258 11452
rect 8314 11450 8338 11452
rect 8394 11450 8418 11452
rect 8474 11450 8498 11452
rect 8554 11450 8560 11452
rect 8314 11398 8316 11450
rect 8496 11398 8498 11450
rect 8252 11396 8258 11398
rect 8314 11396 8338 11398
rect 8394 11396 8418 11398
rect 8474 11396 8498 11398
rect 8554 11396 8560 11398
rect 8252 11387 8560 11396
rect 8864 11354 8892 11698
rect 11173 11452 11481 11461
rect 11173 11450 11179 11452
rect 11235 11450 11259 11452
rect 11315 11450 11339 11452
rect 11395 11450 11419 11452
rect 11475 11450 11481 11452
rect 11235 11398 11237 11450
rect 11417 11398 11419 11450
rect 11173 11396 11179 11398
rect 11235 11396 11259 11398
rect 11315 11396 11339 11398
rect 11395 11396 11419 11398
rect 11475 11396 11481 11398
rect 11173 11387 11481 11396
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 8912 10908 9220 10917
rect 8912 10906 8918 10908
rect 8974 10906 8998 10908
rect 9054 10906 9078 10908
rect 9134 10906 9158 10908
rect 9214 10906 9220 10908
rect 8974 10854 8976 10906
rect 9156 10854 9158 10906
rect 8912 10852 8918 10854
rect 8974 10852 8998 10854
rect 9054 10852 9078 10854
rect 9134 10852 9158 10854
rect 9214 10852 9220 10854
rect 8912 10843 9220 10852
rect 11833 10908 12141 10917
rect 11833 10906 11839 10908
rect 11895 10906 11919 10908
rect 11975 10906 11999 10908
rect 12055 10906 12079 10908
rect 12135 10906 12141 10908
rect 11895 10854 11897 10906
rect 12077 10854 12079 10906
rect 11833 10852 11839 10854
rect 11895 10852 11919 10854
rect 11975 10852 11999 10854
rect 12055 10852 12079 10854
rect 12135 10852 12141 10854
rect 11833 10843 12141 10852
rect 8252 10364 8560 10373
rect 8252 10362 8258 10364
rect 8314 10362 8338 10364
rect 8394 10362 8418 10364
rect 8474 10362 8498 10364
rect 8554 10362 8560 10364
rect 8314 10310 8316 10362
rect 8496 10310 8498 10362
rect 8252 10308 8258 10310
rect 8314 10308 8338 10310
rect 8394 10308 8418 10310
rect 8474 10308 8498 10310
rect 8554 10308 8560 10310
rect 8252 10299 8560 10308
rect 11173 10364 11481 10373
rect 11173 10362 11179 10364
rect 11235 10362 11259 10364
rect 11315 10362 11339 10364
rect 11395 10362 11419 10364
rect 11475 10362 11481 10364
rect 11235 10310 11237 10362
rect 11417 10310 11419 10362
rect 11173 10308 11179 10310
rect 11235 10308 11259 10310
rect 11315 10308 11339 10310
rect 11395 10308 11419 10310
rect 11475 10308 11481 10310
rect 11173 10299 11481 10308
rect 5908 9988 5960 9994
rect 5908 9930 5960 9936
rect 5920 9586 5948 9930
rect 5991 9820 6299 9829
rect 5991 9818 5997 9820
rect 6053 9818 6077 9820
rect 6133 9818 6157 9820
rect 6213 9818 6237 9820
rect 6293 9818 6299 9820
rect 6053 9766 6055 9818
rect 6235 9766 6237 9818
rect 5991 9764 5997 9766
rect 6053 9764 6077 9766
rect 6133 9764 6157 9766
rect 6213 9764 6237 9766
rect 6293 9764 6299 9766
rect 5991 9755 6299 9764
rect 5908 9580 5960 9586
rect 5908 9522 5960 9528
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 5920 8634 5948 9318
rect 6380 8906 6408 9998
rect 6920 9988 6972 9994
rect 8036 9982 8156 10010
rect 6920 9930 6972 9936
rect 6932 9586 6960 9930
rect 7380 9920 7432 9926
rect 7380 9862 7432 9868
rect 8024 9920 8076 9926
rect 8024 9862 8076 9868
rect 7392 9586 7420 9862
rect 8036 9722 8064 9862
rect 8024 9716 8076 9722
rect 8024 9658 8076 9664
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 7208 9178 7236 9454
rect 7472 9376 7524 9382
rect 7472 9318 7524 9324
rect 7484 9178 7512 9318
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7472 9172 7524 9178
rect 7472 9114 7524 9120
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 7196 8968 7248 8974
rect 7196 8910 7248 8916
rect 7932 8968 7984 8974
rect 7932 8910 7984 8916
rect 6368 8900 6420 8906
rect 6368 8842 6420 8848
rect 5991 8732 6299 8741
rect 5991 8730 5997 8732
rect 6053 8730 6077 8732
rect 6133 8730 6157 8732
rect 6213 8730 6237 8732
rect 6293 8730 6299 8732
rect 6053 8678 6055 8730
rect 6235 8678 6237 8730
rect 5991 8676 5997 8678
rect 6053 8676 6077 8678
rect 6133 8676 6157 8678
rect 6213 8676 6237 8678
rect 6293 8676 6299 8678
rect 5991 8667 6299 8676
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 6380 8294 6408 8842
rect 6932 8634 6960 8910
rect 6920 8628 6972 8634
rect 6920 8570 6972 8576
rect 5908 8288 5960 8294
rect 5908 8230 5960 8236
rect 6276 8288 6328 8294
rect 6276 8230 6328 8236
rect 6368 8288 6420 8294
rect 6368 8230 6420 8236
rect 5816 7880 5868 7886
rect 5816 7822 5868 7828
rect 5920 7546 5948 8230
rect 6288 7818 6316 8230
rect 6276 7812 6328 7818
rect 6276 7754 6328 7760
rect 5991 7644 6299 7653
rect 5991 7642 5997 7644
rect 6053 7642 6077 7644
rect 6133 7642 6157 7644
rect 6213 7642 6237 7644
rect 6293 7642 6299 7644
rect 6053 7590 6055 7642
rect 6235 7590 6237 7642
rect 5991 7588 5997 7590
rect 6053 7588 6077 7590
rect 6133 7588 6157 7590
rect 6213 7588 6237 7590
rect 6293 7588 6299 7590
rect 5991 7579 6299 7588
rect 5908 7540 5960 7546
rect 5908 7482 5960 7488
rect 6380 7410 6408 8230
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 6368 7404 6420 7410
rect 6368 7346 6420 7352
rect 6380 7002 6408 7346
rect 6368 6996 6420 7002
rect 6368 6938 6420 6944
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5331 6012 5639 6021
rect 5331 6010 5337 6012
rect 5393 6010 5417 6012
rect 5473 6010 5497 6012
rect 5553 6010 5577 6012
rect 5633 6010 5639 6012
rect 5393 5958 5395 6010
rect 5575 5958 5577 6010
rect 5331 5956 5337 5958
rect 5393 5956 5417 5958
rect 5473 5956 5497 5958
rect 5553 5956 5577 5958
rect 5633 5956 5639 5958
rect 5331 5947 5639 5956
rect 5172 5296 5224 5302
rect 5172 5238 5224 5244
rect 5080 5228 5132 5234
rect 5080 5170 5132 5176
rect 4804 5092 4856 5098
rect 4804 5034 4856 5040
rect 4816 4162 4844 5034
rect 4988 5024 5040 5030
rect 4988 4966 5040 4972
rect 5000 4282 5028 4966
rect 5092 4690 5120 5170
rect 5080 4684 5132 4690
rect 5080 4626 5132 4632
rect 4988 4276 5040 4282
rect 4988 4218 5040 4224
rect 5078 4176 5134 4185
rect 4816 4146 4936 4162
rect 4816 4140 4948 4146
rect 4816 4134 4896 4140
rect 5078 4111 5080 4120
rect 4896 4082 4948 4088
rect 5132 4111 5134 4120
rect 5080 4082 5132 4088
rect 4712 3528 4764 3534
rect 4710 3496 4712 3505
rect 4804 3528 4856 3534
rect 4764 3496 4766 3505
rect 4620 3460 4672 3466
rect 4804 3470 4856 3476
rect 4710 3431 4766 3440
rect 4620 3402 4672 3408
rect 4632 3210 4660 3402
rect 4540 3194 4660 3210
rect 4528 3188 4660 3194
rect 4580 3182 4660 3188
rect 4528 3130 4580 3136
rect 4434 3088 4490 3097
rect 4434 3023 4436 3032
rect 4488 3023 4490 3032
rect 4436 2994 4488 3000
rect 4528 2984 4580 2990
rect 4724 2938 4752 3431
rect 4816 3126 4844 3470
rect 4804 3120 4856 3126
rect 4804 3062 4856 3068
rect 4580 2932 4752 2938
rect 4528 2926 4752 2932
rect 4540 2910 4752 2926
rect 4436 2848 4488 2854
rect 4436 2790 4488 2796
rect 4528 2848 4580 2854
rect 4528 2790 4580 2796
rect 4448 2446 4476 2790
rect 4540 2650 4568 2790
rect 4816 2650 4844 3062
rect 4908 2961 4936 4082
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 5000 3641 5028 3878
rect 4986 3632 5042 3641
rect 4986 3567 5042 3576
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 5000 3126 5028 3334
rect 5092 3194 5120 3878
rect 5184 3534 5212 5238
rect 5331 4924 5639 4933
rect 5331 4922 5337 4924
rect 5393 4922 5417 4924
rect 5473 4922 5497 4924
rect 5553 4922 5577 4924
rect 5633 4922 5639 4924
rect 5393 4870 5395 4922
rect 5575 4870 5577 4922
rect 5331 4868 5337 4870
rect 5393 4868 5417 4870
rect 5473 4868 5497 4870
rect 5553 4868 5577 4870
rect 5633 4868 5639 4870
rect 5331 4859 5639 4868
rect 5736 4826 5764 6598
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 5724 4820 5776 4826
rect 5724 4762 5776 4768
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 5276 4282 5304 4558
rect 5356 4480 5408 4486
rect 5356 4422 5408 4428
rect 5368 4282 5396 4422
rect 5264 4276 5316 4282
rect 5264 4218 5316 4224
rect 5356 4276 5408 4282
rect 5356 4218 5408 4224
rect 5460 4146 5488 4762
rect 5552 4690 5672 4706
rect 5828 4690 5856 6734
rect 5991 6556 6299 6565
rect 5991 6554 5997 6556
rect 6053 6554 6077 6556
rect 6133 6554 6157 6556
rect 6213 6554 6237 6556
rect 6293 6554 6299 6556
rect 6053 6502 6055 6554
rect 6235 6502 6237 6554
rect 5991 6500 5997 6502
rect 6053 6500 6077 6502
rect 6133 6500 6157 6502
rect 6213 6500 6237 6502
rect 6293 6500 6299 6502
rect 5991 6491 6299 6500
rect 7116 6458 7144 7890
rect 7208 7478 7236 8910
rect 7748 8900 7800 8906
rect 7748 8842 7800 8848
rect 7760 7886 7788 8842
rect 7944 8634 7972 8910
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 7748 7880 7800 7886
rect 7748 7822 7800 7828
rect 7656 7812 7708 7818
rect 7656 7754 7708 7760
rect 7196 7472 7248 7478
rect 7196 7414 7248 7420
rect 7288 7200 7340 7206
rect 7288 7142 7340 7148
rect 7300 6798 7328 7142
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 6368 6384 6420 6390
rect 6420 6344 6592 6372
rect 6368 6326 6420 6332
rect 5908 6316 5960 6322
rect 5908 6258 5960 6264
rect 6184 6316 6236 6322
rect 6184 6258 6236 6264
rect 5920 5914 5948 6258
rect 6196 6225 6224 6258
rect 6182 6216 6238 6225
rect 6182 6151 6238 6160
rect 5908 5908 5960 5914
rect 5908 5850 5960 5856
rect 6196 5778 6224 6151
rect 6184 5772 6236 5778
rect 6184 5714 6236 5720
rect 6368 5772 6420 5778
rect 6368 5714 6420 5720
rect 5908 5704 5960 5710
rect 5908 5646 5960 5652
rect 5920 5370 5948 5646
rect 5991 5468 6299 5477
rect 5991 5466 5997 5468
rect 6053 5466 6077 5468
rect 6133 5466 6157 5468
rect 6213 5466 6237 5468
rect 6293 5466 6299 5468
rect 6053 5414 6055 5466
rect 6235 5414 6237 5466
rect 5991 5412 5997 5414
rect 6053 5412 6077 5414
rect 6133 5412 6157 5414
rect 6213 5412 6237 5414
rect 6293 5412 6299 5414
rect 5991 5403 6299 5412
rect 6380 5370 6408 5714
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 5908 5364 5960 5370
rect 5908 5306 5960 5312
rect 6184 5364 6236 5370
rect 6184 5306 6236 5312
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 6092 5160 6144 5166
rect 6092 5102 6144 5108
rect 5540 4684 5672 4690
rect 5592 4678 5672 4684
rect 5540 4626 5592 4632
rect 5540 4548 5592 4554
rect 5540 4490 5592 4496
rect 5552 4282 5580 4490
rect 5644 4298 5672 4678
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 5908 4480 5960 4486
rect 6104 4468 6132 5102
rect 6196 4622 6224 5306
rect 6274 5264 6330 5273
rect 6274 5199 6276 5208
rect 6328 5199 6330 5208
rect 6276 5170 6328 5176
rect 6288 4622 6316 5170
rect 6380 5114 6408 5306
rect 6472 5234 6500 5646
rect 6460 5228 6512 5234
rect 6460 5170 6512 5176
rect 6380 5086 6500 5114
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 5960 4440 6132 4468
rect 5908 4422 5960 4428
rect 5991 4380 6299 4389
rect 5991 4378 5997 4380
rect 6053 4378 6077 4380
rect 6133 4378 6157 4380
rect 6213 4378 6237 4380
rect 6293 4378 6299 4380
rect 6053 4326 6055 4378
rect 6235 4326 6237 4378
rect 5991 4324 5997 4326
rect 6053 4324 6077 4326
rect 6133 4324 6157 4326
rect 6213 4324 6237 4326
rect 6293 4324 6299 4326
rect 5991 4315 6299 4324
rect 5540 4276 5592 4282
rect 5644 4270 5856 4298
rect 5540 4218 5592 4224
rect 5722 4176 5778 4185
rect 5644 4146 5722 4162
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5632 4140 5722 4146
rect 5684 4134 5722 4140
rect 5722 4111 5778 4120
rect 5632 4082 5684 4088
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 5331 3836 5639 3845
rect 5331 3834 5337 3836
rect 5393 3834 5417 3836
rect 5473 3834 5497 3836
rect 5553 3834 5577 3836
rect 5633 3834 5639 3836
rect 5393 3782 5395 3834
rect 5575 3782 5577 3834
rect 5331 3780 5337 3782
rect 5393 3780 5417 3782
rect 5473 3780 5497 3782
rect 5553 3780 5577 3782
rect 5633 3780 5639 3782
rect 5331 3771 5639 3780
rect 5736 3738 5764 3878
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5172 3528 5224 3534
rect 5172 3470 5224 3476
rect 5724 3460 5776 3466
rect 5724 3402 5776 3408
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 4988 3120 5040 3126
rect 4988 3062 5040 3068
rect 5736 3058 5764 3402
rect 5080 3052 5132 3058
rect 5080 2994 5132 3000
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 4988 2984 5040 2990
rect 4894 2952 4950 2961
rect 4988 2926 5040 2932
rect 4894 2887 4950 2896
rect 4528 2644 4580 2650
rect 4528 2586 4580 2592
rect 4804 2644 4856 2650
rect 4804 2586 4856 2592
rect 4436 2440 4488 2446
rect 4436 2382 4488 2388
rect 5000 2378 5028 2926
rect 5092 2825 5120 2994
rect 5078 2816 5134 2825
rect 5078 2751 5134 2760
rect 5331 2748 5639 2757
rect 5331 2746 5337 2748
rect 5393 2746 5417 2748
rect 5473 2746 5497 2748
rect 5553 2746 5577 2748
rect 5633 2746 5639 2748
rect 5393 2694 5395 2746
rect 5575 2694 5577 2746
rect 5331 2692 5337 2694
rect 5393 2692 5417 2694
rect 5473 2692 5497 2694
rect 5553 2692 5577 2694
rect 5633 2692 5639 2694
rect 5331 2683 5639 2692
rect 5448 2576 5500 2582
rect 5448 2518 5500 2524
rect 5460 2378 5488 2518
rect 5736 2446 5764 2994
rect 5828 2990 5856 4270
rect 6380 4078 6408 4966
rect 6472 4826 6500 5086
rect 6460 4820 6512 4826
rect 6460 4762 6512 4768
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 6368 4072 6420 4078
rect 6368 4014 6420 4020
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 6276 3936 6328 3942
rect 6276 3878 6328 3884
rect 5908 3664 5960 3670
rect 5908 3606 5960 3612
rect 5920 3126 5948 3606
rect 6104 3534 6132 3878
rect 6092 3528 6144 3534
rect 6092 3470 6144 3476
rect 6288 3380 6316 3878
rect 6288 3352 6408 3380
rect 5991 3292 6299 3301
rect 5991 3290 5997 3292
rect 6053 3290 6077 3292
rect 6133 3290 6157 3292
rect 6213 3290 6237 3292
rect 6293 3290 6299 3292
rect 6053 3238 6055 3290
rect 6235 3238 6237 3290
rect 5991 3236 5997 3238
rect 6053 3236 6077 3238
rect 6133 3236 6157 3238
rect 6213 3236 6237 3238
rect 6293 3236 6299 3238
rect 5991 3227 6299 3236
rect 6380 3194 6408 3352
rect 6368 3188 6420 3194
rect 6368 3130 6420 3136
rect 5908 3120 5960 3126
rect 5908 3062 5960 3068
rect 6472 3058 6500 4082
rect 6564 4026 6592 6344
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 6644 6248 6696 6254
rect 7576 6225 7604 6258
rect 6644 6190 6696 6196
rect 7562 6216 7618 6225
rect 6656 5914 6684 6190
rect 7562 6151 7618 6160
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 6656 5710 6684 5850
rect 6920 5840 6972 5846
rect 6920 5782 6972 5788
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6748 5302 6776 5510
rect 6932 5370 6960 5782
rect 7104 5704 7156 5710
rect 7104 5646 7156 5652
rect 7288 5704 7340 5710
rect 7288 5646 7340 5652
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 6736 5296 6788 5302
rect 6736 5238 6788 5244
rect 6918 5264 6974 5273
rect 6918 5199 6920 5208
rect 6972 5199 6974 5208
rect 6920 5170 6972 5176
rect 6644 5024 6696 5030
rect 6644 4966 6696 4972
rect 6656 4690 6684 4966
rect 6644 4684 6696 4690
rect 6644 4626 6696 4632
rect 6828 4548 6880 4554
rect 6828 4490 6880 4496
rect 6840 4214 6868 4490
rect 6828 4208 6880 4214
rect 6828 4150 6880 4156
rect 6564 3998 6684 4026
rect 6552 3732 6604 3738
rect 6552 3674 6604 3680
rect 6564 3194 6592 3674
rect 6656 3194 6684 3998
rect 6736 3936 6788 3942
rect 6932 3924 6960 5170
rect 7116 5137 7144 5646
rect 7102 5128 7158 5137
rect 7300 5098 7328 5646
rect 7102 5063 7104 5072
rect 7156 5063 7158 5072
rect 7288 5092 7340 5098
rect 7104 5034 7156 5040
rect 7288 5034 7340 5040
rect 7116 4214 7144 5034
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7484 4622 7512 4966
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 7576 4486 7604 6151
rect 7668 5710 7696 7754
rect 7760 7410 7788 7822
rect 7852 7546 7880 8434
rect 8128 7886 8156 9982
rect 8912 9820 9220 9829
rect 8912 9818 8918 9820
rect 8974 9818 8998 9820
rect 9054 9818 9078 9820
rect 9134 9818 9158 9820
rect 9214 9818 9220 9820
rect 8974 9766 8976 9818
rect 9156 9766 9158 9818
rect 8912 9764 8918 9766
rect 8974 9764 8998 9766
rect 9054 9764 9078 9766
rect 9134 9764 9158 9766
rect 9214 9764 9220 9766
rect 8912 9755 9220 9764
rect 11833 9820 12141 9829
rect 11833 9818 11839 9820
rect 11895 9818 11919 9820
rect 11975 9818 11999 9820
rect 12055 9818 12079 9820
rect 12135 9818 12141 9820
rect 11895 9766 11897 9818
rect 12077 9766 12079 9818
rect 11833 9764 11839 9766
rect 11895 9764 11919 9766
rect 11975 9764 11999 9766
rect 12055 9764 12079 9766
rect 12135 9764 12141 9766
rect 11833 9755 12141 9764
rect 8252 9276 8560 9285
rect 8252 9274 8258 9276
rect 8314 9274 8338 9276
rect 8394 9274 8418 9276
rect 8474 9274 8498 9276
rect 8554 9274 8560 9276
rect 8314 9222 8316 9274
rect 8496 9222 8498 9274
rect 8252 9220 8258 9222
rect 8314 9220 8338 9222
rect 8394 9220 8418 9222
rect 8474 9220 8498 9222
rect 8554 9220 8560 9222
rect 8252 9211 8560 9220
rect 11173 9276 11481 9285
rect 11173 9274 11179 9276
rect 11235 9274 11259 9276
rect 11315 9274 11339 9276
rect 11395 9274 11419 9276
rect 11475 9274 11481 9276
rect 11235 9222 11237 9274
rect 11417 9222 11419 9274
rect 11173 9220 11179 9222
rect 11235 9220 11259 9222
rect 11315 9220 11339 9222
rect 11395 9220 11419 9222
rect 11475 9220 11481 9222
rect 11173 9211 11481 9220
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 9312 8968 9364 8974
rect 9312 8910 9364 8916
rect 8772 8634 8800 8910
rect 8912 8732 9220 8741
rect 8912 8730 8918 8732
rect 8974 8730 8998 8732
rect 9054 8730 9078 8732
rect 9134 8730 9158 8732
rect 9214 8730 9220 8732
rect 8974 8678 8976 8730
rect 9156 8678 9158 8730
rect 8912 8676 8918 8678
rect 8974 8676 8998 8678
rect 9054 8676 9078 8678
rect 9134 8676 9158 8678
rect 9214 8676 9220 8678
rect 8912 8667 9220 8676
rect 8760 8628 8812 8634
rect 8760 8570 8812 8576
rect 8576 8288 8628 8294
rect 8576 8230 8628 8236
rect 8252 8188 8560 8197
rect 8252 8186 8258 8188
rect 8314 8186 8338 8188
rect 8394 8186 8418 8188
rect 8474 8186 8498 8188
rect 8554 8186 8560 8188
rect 8314 8134 8316 8186
rect 8496 8134 8498 8186
rect 8252 8132 8258 8134
rect 8314 8132 8338 8134
rect 8394 8132 8418 8134
rect 8474 8132 8498 8134
rect 8554 8132 8560 8134
rect 8252 8123 8560 8132
rect 8588 7954 8616 8230
rect 8576 7948 8628 7954
rect 8576 7890 8628 7896
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 7840 7540 7892 7546
rect 7840 7482 7892 7488
rect 8128 7426 8156 7822
rect 9324 7818 9352 8910
rect 9956 8900 10008 8906
rect 9956 8842 10008 8848
rect 9968 8634 9996 8842
rect 11833 8732 12141 8741
rect 11833 8730 11839 8732
rect 11895 8730 11919 8732
rect 11975 8730 11999 8732
rect 12055 8730 12079 8732
rect 12135 8730 12141 8732
rect 11895 8678 11897 8730
rect 12077 8678 12079 8730
rect 11833 8676 11839 8678
rect 11895 8676 11919 8678
rect 11975 8676 11999 8678
rect 12055 8676 12079 8678
rect 12135 8676 12141 8678
rect 11833 8667 12141 8676
rect 9956 8628 10008 8634
rect 9956 8570 10008 8576
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 10060 8090 10088 8434
rect 11173 8188 11481 8197
rect 11173 8186 11179 8188
rect 11235 8186 11259 8188
rect 11315 8186 11339 8188
rect 11395 8186 11419 8188
rect 11475 8186 11481 8188
rect 11235 8134 11237 8186
rect 11417 8134 11419 8186
rect 11173 8132 11179 8134
rect 11235 8132 11259 8134
rect 11315 8132 11339 8134
rect 11395 8132 11419 8134
rect 11475 8132 11481 8134
rect 11173 8123 11481 8132
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 9312 7812 9364 7818
rect 9312 7754 9364 7760
rect 8912 7644 9220 7653
rect 8912 7642 8918 7644
rect 8974 7642 8998 7644
rect 9054 7642 9078 7644
rect 9134 7642 9158 7644
rect 9214 7642 9220 7644
rect 8974 7590 8976 7642
rect 9156 7590 9158 7642
rect 8912 7588 8918 7590
rect 8974 7588 8998 7590
rect 9054 7588 9078 7590
rect 9134 7588 9158 7590
rect 9214 7588 9220 7590
rect 8912 7579 9220 7588
rect 11833 7644 12141 7653
rect 11833 7642 11839 7644
rect 11895 7642 11919 7644
rect 11975 7642 11999 7644
rect 12055 7642 12079 7644
rect 12135 7642 12141 7644
rect 11895 7590 11897 7642
rect 12077 7590 12079 7642
rect 11833 7588 11839 7590
rect 11895 7588 11919 7590
rect 11975 7588 11999 7590
rect 12055 7588 12079 7590
rect 12135 7588 12141 7590
rect 11833 7579 12141 7588
rect 8036 7410 8156 7426
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 8024 7404 8156 7410
rect 8076 7398 8156 7404
rect 8852 7404 8904 7410
rect 8024 7346 8076 7352
rect 8852 7346 8904 7352
rect 9588 7404 9640 7410
rect 9588 7346 9640 7352
rect 11060 7404 11112 7410
rect 11060 7346 11112 7352
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 8760 7336 8812 7342
rect 8760 7278 8812 7284
rect 8252 7100 8560 7109
rect 8252 7098 8258 7100
rect 8314 7098 8338 7100
rect 8394 7098 8418 7100
rect 8474 7098 8498 7100
rect 8554 7098 8560 7100
rect 8314 7046 8316 7098
rect 8496 7046 8498 7098
rect 8252 7044 8258 7046
rect 8314 7044 8338 7046
rect 8394 7044 8418 7046
rect 8474 7044 8498 7046
rect 8554 7044 8560 7046
rect 8252 7035 8560 7044
rect 7840 6452 7892 6458
rect 7840 6394 7892 6400
rect 7656 5704 7708 5710
rect 7748 5704 7800 5710
rect 7656 5646 7708 5652
rect 7746 5672 7748 5681
rect 7800 5672 7802 5681
rect 7668 5216 7696 5646
rect 7746 5607 7802 5616
rect 7760 5574 7788 5607
rect 7852 5574 7880 6394
rect 8588 6361 8616 7278
rect 8680 7002 8708 7278
rect 8668 6996 8720 7002
rect 8668 6938 8720 6944
rect 8772 6934 8800 7278
rect 8760 6928 8812 6934
rect 8760 6870 8812 6876
rect 8668 6656 8720 6662
rect 8668 6598 8720 6604
rect 8574 6352 8630 6361
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 8116 6316 8168 6322
rect 8574 6287 8630 6296
rect 8116 6258 8168 6264
rect 7932 6112 7984 6118
rect 7932 6054 7984 6060
rect 7748 5568 7800 5574
rect 7748 5510 7800 5516
rect 7840 5568 7892 5574
rect 7840 5510 7892 5516
rect 7852 5370 7880 5510
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 7852 5234 7880 5306
rect 7748 5228 7800 5234
rect 7668 5188 7748 5216
rect 7668 4622 7696 5188
rect 7748 5170 7800 5176
rect 7840 5228 7892 5234
rect 7840 5170 7892 5176
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 7656 4616 7708 4622
rect 7656 4558 7708 4564
rect 7564 4480 7616 4486
rect 7564 4422 7616 4428
rect 7760 4282 7788 4966
rect 7852 4622 7880 5170
rect 7840 4616 7892 4622
rect 7840 4558 7892 4564
rect 7748 4276 7800 4282
rect 7748 4218 7800 4224
rect 7104 4208 7156 4214
rect 7104 4150 7156 4156
rect 7012 3936 7064 3942
rect 6932 3896 7012 3924
rect 6736 3878 6788 3884
rect 7012 3878 7064 3884
rect 7656 3936 7708 3942
rect 7656 3878 7708 3884
rect 6748 3602 6776 3878
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 7010 3632 7066 3641
rect 6736 3596 6788 3602
rect 7010 3567 7066 3576
rect 6736 3538 6788 3544
rect 6552 3188 6604 3194
rect 6552 3130 6604 3136
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 6656 3058 6684 3130
rect 6092 3052 6144 3058
rect 6092 2994 6144 3000
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 5816 2984 5868 2990
rect 5816 2926 5868 2932
rect 5828 2854 5856 2926
rect 6000 2916 6052 2922
rect 6000 2858 6052 2864
rect 5816 2848 5868 2854
rect 5816 2790 5868 2796
rect 6012 2446 6040 2858
rect 6104 2582 6132 2994
rect 6092 2576 6144 2582
rect 6092 2518 6144 2524
rect 6748 2514 6776 3538
rect 7024 2922 7052 3567
rect 7300 3126 7328 3674
rect 7472 3664 7524 3670
rect 7472 3606 7524 3612
rect 7484 3534 7512 3606
rect 7668 3534 7696 3878
rect 7760 3738 7788 4218
rect 7944 4214 7972 6054
rect 8036 5574 8064 6258
rect 8128 5914 8156 6258
rect 8208 6248 8260 6254
rect 8260 6196 8616 6202
rect 8208 6190 8616 6196
rect 8220 6174 8616 6190
rect 8252 6012 8560 6021
rect 8252 6010 8258 6012
rect 8314 6010 8338 6012
rect 8394 6010 8418 6012
rect 8474 6010 8498 6012
rect 8554 6010 8560 6012
rect 8314 5958 8316 6010
rect 8496 5958 8498 6010
rect 8252 5956 8258 5958
rect 8314 5956 8338 5958
rect 8394 5956 8418 5958
rect 8474 5956 8498 5958
rect 8554 5956 8560 5958
rect 8252 5947 8560 5956
rect 8116 5908 8168 5914
rect 8116 5850 8168 5856
rect 8392 5772 8444 5778
rect 8392 5714 8444 5720
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 8024 5568 8076 5574
rect 8024 5510 8076 5516
rect 8128 4978 8156 5646
rect 8404 5137 8432 5714
rect 8588 5234 8616 6174
rect 8680 5710 8708 6598
rect 8772 5778 8800 6870
rect 8864 6730 8892 7346
rect 9600 6798 9628 7346
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 8852 6724 8904 6730
rect 8852 6666 8904 6672
rect 9312 6724 9364 6730
rect 9312 6666 9364 6672
rect 8912 6556 9220 6565
rect 8912 6554 8918 6556
rect 8974 6554 8998 6556
rect 9054 6554 9078 6556
rect 9134 6554 9158 6556
rect 9214 6554 9220 6556
rect 8974 6502 8976 6554
rect 9156 6502 9158 6554
rect 8912 6500 8918 6502
rect 8974 6500 8998 6502
rect 9054 6500 9078 6502
rect 9134 6500 9158 6502
rect 9214 6500 9220 6502
rect 8912 6491 9220 6500
rect 9034 6352 9090 6361
rect 8852 6316 8904 6322
rect 9324 6322 9352 6666
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 9034 6287 9036 6296
rect 8852 6258 8904 6264
rect 9088 6287 9090 6296
rect 9312 6316 9364 6322
rect 9036 6258 9088 6264
rect 9312 6258 9364 6264
rect 8864 5846 8892 6258
rect 8942 6216 8998 6225
rect 8942 6151 8998 6160
rect 9312 6180 9364 6186
rect 8956 6118 8984 6151
rect 9312 6122 9364 6128
rect 8944 6112 8996 6118
rect 8944 6054 8996 6060
rect 8852 5840 8904 5846
rect 8852 5782 8904 5788
rect 8760 5772 8812 5778
rect 8760 5714 8812 5720
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 8576 5228 8628 5234
rect 8576 5170 8628 5176
rect 8390 5128 8446 5137
rect 8390 5063 8446 5072
rect 8404 5030 8432 5063
rect 8036 4950 8156 4978
rect 8392 5024 8444 5030
rect 8392 4966 8444 4972
rect 8036 4554 8064 4950
rect 8252 4924 8560 4933
rect 8252 4922 8258 4924
rect 8314 4922 8338 4924
rect 8394 4922 8418 4924
rect 8474 4922 8498 4924
rect 8554 4922 8560 4924
rect 8314 4870 8316 4922
rect 8496 4870 8498 4922
rect 8252 4868 8258 4870
rect 8314 4868 8338 4870
rect 8394 4868 8418 4870
rect 8474 4868 8498 4870
rect 8554 4868 8560 4870
rect 8252 4859 8560 4868
rect 8116 4752 8168 4758
rect 8116 4694 8168 4700
rect 8024 4548 8076 4554
rect 8024 4490 8076 4496
rect 7932 4208 7984 4214
rect 7930 4176 7932 4185
rect 7984 4176 7986 4185
rect 7930 4111 7986 4120
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 8128 3670 8156 4694
rect 8484 4616 8536 4622
rect 8484 4558 8536 4564
rect 8496 4214 8524 4558
rect 8484 4208 8536 4214
rect 8484 4150 8536 4156
rect 8252 3836 8560 3845
rect 8252 3834 8258 3836
rect 8314 3834 8338 3836
rect 8394 3834 8418 3836
rect 8474 3834 8498 3836
rect 8554 3834 8560 3836
rect 8314 3782 8316 3834
rect 8496 3782 8498 3834
rect 8252 3780 8258 3782
rect 8314 3780 8338 3782
rect 8394 3780 8418 3782
rect 8474 3780 8498 3782
rect 8554 3780 8560 3782
rect 8252 3771 8560 3780
rect 8116 3664 8168 3670
rect 8116 3606 8168 3612
rect 8588 3534 8616 5170
rect 8668 4480 8720 4486
rect 8668 4422 8720 4428
rect 8680 4146 8708 4422
rect 8772 4162 8800 5714
rect 9324 5681 9352 6122
rect 9310 5672 9366 5681
rect 9310 5607 9366 5616
rect 8912 5468 9220 5477
rect 8912 5466 8918 5468
rect 8974 5466 8998 5468
rect 9054 5466 9078 5468
rect 9134 5466 9158 5468
rect 9214 5466 9220 5468
rect 8974 5414 8976 5466
rect 9156 5414 9158 5466
rect 8912 5412 8918 5414
rect 8974 5412 8998 5414
rect 9054 5412 9078 5414
rect 9134 5412 9158 5414
rect 9214 5412 9220 5414
rect 8912 5403 9220 5412
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 9220 5228 9272 5234
rect 9220 5170 9272 5176
rect 8956 4758 8984 5170
rect 8944 4752 8996 4758
rect 8944 4694 8996 4700
rect 8956 4593 8984 4694
rect 9232 4690 9260 5170
rect 9324 4826 9352 5607
rect 9312 4820 9364 4826
rect 9312 4762 9364 4768
rect 9220 4684 9272 4690
rect 9220 4626 9272 4632
rect 8942 4584 8998 4593
rect 8942 4519 8998 4528
rect 8912 4380 9220 4389
rect 8912 4378 8918 4380
rect 8974 4378 8998 4380
rect 9054 4378 9078 4380
rect 9134 4378 9158 4380
rect 9214 4378 9220 4380
rect 8974 4326 8976 4378
rect 9156 4326 9158 4378
rect 8912 4324 8918 4326
rect 8974 4324 8998 4326
rect 9054 4324 9078 4326
rect 9134 4324 9158 4326
rect 9214 4324 9220 4326
rect 8912 4315 9220 4324
rect 8944 4276 8996 4282
rect 8944 4218 8996 4224
rect 8772 4146 8892 4162
rect 8668 4140 8720 4146
rect 8668 4082 8720 4088
rect 8772 4140 8904 4146
rect 8772 4134 8852 4140
rect 8668 3936 8720 3942
rect 8668 3878 8720 3884
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7656 3528 7708 3534
rect 7932 3528 7984 3534
rect 7656 3470 7708 3476
rect 7930 3496 7932 3505
rect 8576 3528 8628 3534
rect 7984 3496 7986 3505
rect 7484 3126 7512 3470
rect 7986 3454 8156 3482
rect 8576 3470 8628 3476
rect 7930 3431 7986 3440
rect 7932 3392 7984 3398
rect 7932 3334 7984 3340
rect 7944 3194 7972 3334
rect 7932 3188 7984 3194
rect 7932 3130 7984 3136
rect 7288 3120 7340 3126
rect 7288 3062 7340 3068
rect 7472 3120 7524 3126
rect 7472 3062 7524 3068
rect 7012 2916 7064 2922
rect 7012 2858 7064 2864
rect 6920 2848 6972 2854
rect 6972 2796 7052 2802
rect 6920 2790 7052 2796
rect 6932 2774 7052 2790
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 7024 2446 7052 2774
rect 8128 2650 8156 3454
rect 8576 2984 8628 2990
rect 8576 2926 8628 2932
rect 8252 2748 8560 2757
rect 8252 2746 8258 2748
rect 8314 2746 8338 2748
rect 8394 2746 8418 2748
rect 8474 2746 8498 2748
rect 8554 2746 8560 2748
rect 8314 2694 8316 2746
rect 8496 2694 8498 2746
rect 8252 2692 8258 2694
rect 8314 2692 8338 2694
rect 8394 2692 8418 2694
rect 8474 2692 8498 2694
rect 8554 2692 8560 2694
rect 8252 2683 8560 2692
rect 8588 2650 8616 2926
rect 8680 2650 8708 3878
rect 8772 3602 8800 4134
rect 8852 4082 8904 4088
rect 8760 3596 8812 3602
rect 8760 3538 8812 3544
rect 8772 3058 8800 3538
rect 8956 3398 8984 4218
rect 9324 4214 9352 4762
rect 9416 4486 9444 6598
rect 9634 6384 9686 6390
rect 9686 6332 9720 6338
rect 9634 6326 9720 6332
rect 9646 6310 9720 6326
rect 9496 6248 9548 6254
rect 9692 6225 9720 6310
rect 9496 6190 9548 6196
rect 9678 6216 9734 6225
rect 9508 5370 9536 6190
rect 9678 6151 9734 6160
rect 9588 5636 9640 5642
rect 9588 5578 9640 5584
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 9600 5234 9628 5578
rect 9588 5228 9640 5234
rect 9588 5170 9640 5176
rect 9496 5024 9548 5030
rect 9496 4966 9548 4972
rect 9508 4826 9536 4966
rect 9496 4820 9548 4826
rect 9496 4762 9548 4768
rect 9600 4672 9628 5170
rect 9784 5166 9812 7142
rect 9956 6928 10008 6934
rect 9956 6870 10008 6876
rect 9864 6384 9916 6390
rect 9864 6326 9916 6332
rect 9876 6254 9904 6326
rect 9864 6248 9916 6254
rect 9864 6190 9916 6196
rect 9968 5574 9996 6870
rect 11072 6798 11100 7346
rect 11173 7100 11481 7109
rect 11173 7098 11179 7100
rect 11235 7098 11259 7100
rect 11315 7098 11339 7100
rect 11395 7098 11419 7100
rect 11475 7098 11481 7100
rect 11235 7046 11237 7098
rect 11417 7046 11419 7098
rect 11173 7044 11179 7046
rect 11235 7044 11259 7046
rect 11315 7044 11339 7046
rect 11395 7044 11419 7046
rect 11475 7044 11481 7046
rect 11173 7035 11481 7044
rect 12268 6866 12296 13126
rect 12256 6860 12308 6866
rect 12256 6802 12308 6808
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 11833 6556 12141 6565
rect 11833 6554 11839 6556
rect 11895 6554 11919 6556
rect 11975 6554 11999 6556
rect 12055 6554 12079 6556
rect 12135 6554 12141 6556
rect 11895 6502 11897 6554
rect 12077 6502 12079 6554
rect 11833 6500 11839 6502
rect 11895 6500 11919 6502
rect 11975 6500 11999 6502
rect 12055 6500 12079 6502
rect 12135 6500 12141 6502
rect 11833 6491 12141 6500
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 9864 5568 9916 5574
rect 9864 5510 9916 5516
rect 9956 5568 10008 5574
rect 9956 5510 10008 5516
rect 9772 5160 9824 5166
rect 9772 5102 9824 5108
rect 9876 4826 9904 5510
rect 9968 5166 9996 5510
rect 9956 5160 10008 5166
rect 9956 5102 10008 5108
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9864 4820 9916 4826
rect 9864 4762 9916 4768
rect 9508 4644 9628 4672
rect 9680 4684 9732 4690
rect 9404 4480 9456 4486
rect 9404 4422 9456 4428
rect 9402 4312 9458 4321
rect 9508 4282 9536 4644
rect 9680 4626 9732 4632
rect 9588 4548 9640 4554
rect 9588 4490 9640 4496
rect 9402 4247 9458 4256
rect 9496 4276 9548 4282
rect 9312 4208 9364 4214
rect 9312 4150 9364 4156
rect 9036 4140 9088 4146
rect 9036 4082 9088 4088
rect 9048 3466 9076 4082
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 9036 3460 9088 3466
rect 9036 3402 9088 3408
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 8912 3292 9220 3301
rect 8912 3290 8918 3292
rect 8974 3290 8998 3292
rect 9054 3290 9078 3292
rect 9134 3290 9158 3292
rect 9214 3290 9220 3292
rect 8974 3238 8976 3290
rect 9156 3238 9158 3290
rect 8912 3236 8918 3238
rect 8974 3236 8998 3238
rect 9054 3236 9078 3238
rect 9134 3236 9158 3238
rect 9214 3236 9220 3238
rect 8912 3227 9220 3236
rect 8760 3052 8812 3058
rect 8760 2994 8812 3000
rect 9034 2952 9090 2961
rect 9034 2887 9090 2896
rect 9048 2650 9076 2887
rect 8116 2644 8168 2650
rect 8116 2586 8168 2592
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 9324 2446 9352 3470
rect 9416 2514 9444 4247
rect 9496 4218 9548 4224
rect 9508 3602 9536 4218
rect 9600 3738 9628 4490
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9496 3596 9548 3602
rect 9496 3538 9548 3544
rect 9496 3392 9548 3398
rect 9496 3334 9548 3340
rect 9508 3194 9536 3334
rect 9496 3188 9548 3194
rect 9496 3130 9548 3136
rect 9404 2508 9456 2514
rect 9404 2450 9456 2456
rect 9600 2446 9628 3674
rect 9692 2922 9720 4626
rect 9680 2916 9732 2922
rect 9680 2858 9732 2864
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 6000 2440 6052 2446
rect 6000 2382 6052 2388
rect 7012 2440 7064 2446
rect 7012 2382 7064 2388
rect 9312 2440 9364 2446
rect 9312 2382 9364 2388
rect 9588 2440 9640 2446
rect 9588 2382 9640 2388
rect 4988 2372 5040 2378
rect 4988 2314 5040 2320
rect 5448 2372 5500 2378
rect 5448 2314 5500 2320
rect 5460 2038 5488 2314
rect 5828 2106 5856 2382
rect 9784 2310 9812 4762
rect 10060 4622 10088 6394
rect 10232 6248 10284 6254
rect 10230 6216 10232 6225
rect 10284 6216 10286 6225
rect 10230 6151 10286 6160
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 11072 5914 11100 6054
rect 11173 6012 11481 6021
rect 11173 6010 11179 6012
rect 11235 6010 11259 6012
rect 11315 6010 11339 6012
rect 11395 6010 11419 6012
rect 11475 6010 11481 6012
rect 11235 5958 11237 6010
rect 11417 5958 11419 6010
rect 11173 5956 11179 5958
rect 11235 5956 11259 5958
rect 11315 5956 11339 5958
rect 11395 5956 11419 5958
rect 11475 5956 11481 5958
rect 11173 5947 11481 5956
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 10508 5772 10560 5778
rect 10508 5714 10560 5720
rect 10324 5704 10376 5710
rect 10520 5658 10548 5714
rect 10324 5646 10376 5652
rect 10336 5574 10364 5646
rect 10428 5630 10548 5658
rect 10428 5574 10456 5630
rect 10324 5568 10376 5574
rect 10324 5510 10376 5516
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 10508 5568 10560 5574
rect 10508 5510 10560 5516
rect 10428 5234 10456 5510
rect 10520 5370 10548 5510
rect 11833 5468 12141 5477
rect 11833 5466 11839 5468
rect 11895 5466 11919 5468
rect 11975 5466 11999 5468
rect 12055 5466 12079 5468
rect 12135 5466 12141 5468
rect 11895 5414 11897 5466
rect 12077 5414 12079 5466
rect 11833 5412 11839 5414
rect 11895 5412 11919 5414
rect 11975 5412 11999 5414
rect 12055 5412 12079 5414
rect 12135 5412 12141 5414
rect 11833 5403 12141 5412
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10416 5228 10468 5234
rect 10416 5170 10468 5176
rect 11173 4924 11481 4933
rect 11173 4922 11179 4924
rect 11235 4922 11259 4924
rect 11315 4922 11339 4924
rect 11395 4922 11419 4924
rect 11475 4922 11481 4924
rect 11235 4870 11237 4922
rect 11417 4870 11419 4922
rect 11173 4868 11179 4870
rect 11235 4868 11259 4870
rect 11315 4868 11339 4870
rect 11395 4868 11419 4870
rect 11475 4868 11481 4870
rect 11173 4859 11481 4868
rect 10048 4616 10100 4622
rect 10048 4558 10100 4564
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 10048 4480 10100 4486
rect 10048 4422 10100 4428
rect 10060 4214 10088 4422
rect 10048 4208 10100 4214
rect 10048 4150 10100 4156
rect 10244 3738 10272 4558
rect 11833 4380 12141 4389
rect 11833 4378 11839 4380
rect 11895 4378 11919 4380
rect 11975 4378 11999 4380
rect 12055 4378 12079 4380
rect 12135 4378 12141 4380
rect 11895 4326 11897 4378
rect 12077 4326 12079 4378
rect 11833 4324 11839 4326
rect 11895 4324 11919 4326
rect 11975 4324 11999 4326
rect 12055 4324 12079 4326
rect 12135 4324 12141 4326
rect 11833 4315 12141 4324
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10232 3732 10284 3738
rect 10232 3674 10284 3680
rect 10612 3466 10640 3878
rect 11173 3836 11481 3845
rect 11173 3834 11179 3836
rect 11235 3834 11259 3836
rect 11315 3834 11339 3836
rect 11395 3834 11419 3836
rect 11475 3834 11481 3836
rect 11235 3782 11237 3834
rect 11417 3782 11419 3834
rect 11173 3780 11179 3782
rect 11235 3780 11259 3782
rect 11315 3780 11339 3782
rect 11395 3780 11419 3782
rect 11475 3780 11481 3782
rect 11173 3771 11481 3780
rect 12256 3528 12308 3534
rect 12256 3470 12308 3476
rect 10600 3460 10652 3466
rect 10600 3402 10652 3408
rect 11833 3292 12141 3301
rect 11833 3290 11839 3292
rect 11895 3290 11919 3292
rect 11975 3290 11999 3292
rect 12055 3290 12079 3292
rect 12135 3290 12141 3292
rect 11895 3238 11897 3290
rect 12077 3238 12079 3290
rect 11833 3236 11839 3238
rect 11895 3236 11919 3238
rect 11975 3236 11999 3238
rect 12055 3236 12079 3238
rect 12135 3236 12141 3238
rect 11833 3227 12141 3236
rect 11173 2748 11481 2757
rect 11173 2746 11179 2748
rect 11235 2746 11259 2748
rect 11315 2746 11339 2748
rect 11395 2746 11419 2748
rect 11475 2746 11481 2748
rect 11235 2694 11237 2746
rect 11417 2694 11419 2746
rect 11173 2692 11179 2694
rect 11235 2692 11259 2694
rect 11315 2692 11339 2694
rect 11395 2692 11419 2694
rect 11475 2692 11481 2694
rect 11173 2683 11481 2692
rect 12268 2650 12296 3470
rect 12256 2644 12308 2650
rect 12256 2586 12308 2592
rect 9772 2304 9824 2310
rect 9772 2246 9824 2252
rect 12808 2304 12860 2310
rect 12808 2246 12860 2252
rect 5991 2204 6299 2213
rect 5991 2202 5997 2204
rect 6053 2202 6077 2204
rect 6133 2202 6157 2204
rect 6213 2202 6237 2204
rect 6293 2202 6299 2204
rect 6053 2150 6055 2202
rect 6235 2150 6237 2202
rect 5991 2148 5997 2150
rect 6053 2148 6077 2150
rect 6133 2148 6157 2150
rect 6213 2148 6237 2150
rect 6293 2148 6299 2150
rect 5991 2139 6299 2148
rect 8912 2204 9220 2213
rect 8912 2202 8918 2204
rect 8974 2202 8998 2204
rect 9054 2202 9078 2204
rect 9134 2202 9158 2204
rect 9214 2202 9220 2204
rect 8974 2150 8976 2202
rect 9156 2150 9158 2202
rect 8912 2148 8918 2150
rect 8974 2148 8998 2150
rect 9054 2148 9078 2150
rect 9134 2148 9158 2150
rect 9214 2148 9220 2150
rect 8912 2139 9220 2148
rect 11833 2204 12141 2213
rect 11833 2202 11839 2204
rect 11895 2202 11919 2204
rect 11975 2202 11999 2204
rect 12055 2202 12079 2204
rect 12135 2202 12141 2204
rect 11895 2150 11897 2202
rect 12077 2150 12079 2202
rect 11833 2148 11839 2150
rect 11895 2148 11919 2150
rect 11975 2148 11999 2150
rect 12055 2148 12079 2150
rect 12135 2148 12141 2150
rect 11833 2139 12141 2148
rect 5816 2100 5868 2106
rect 5816 2042 5868 2048
rect 4344 2032 4396 2038
rect 4344 1974 4396 1980
rect 5448 2032 5500 2038
rect 5448 1974 5500 1980
rect 18 0 74 800
rect 12820 785 12848 2246
rect 12806 776 12862 785
rect 12806 711 12862 720
<< via2 >>
rect 4066 15000 4122 15056
rect 2416 13626 2472 13628
rect 2496 13626 2552 13628
rect 2576 13626 2632 13628
rect 2656 13626 2712 13628
rect 2416 13574 2462 13626
rect 2462 13574 2472 13626
rect 2496 13574 2526 13626
rect 2526 13574 2538 13626
rect 2538 13574 2552 13626
rect 2576 13574 2590 13626
rect 2590 13574 2602 13626
rect 2602 13574 2632 13626
rect 2656 13574 2666 13626
rect 2666 13574 2712 13626
rect 2416 13572 2472 13574
rect 2496 13572 2552 13574
rect 2576 13572 2632 13574
rect 2656 13572 2712 13574
rect 5337 13626 5393 13628
rect 5417 13626 5473 13628
rect 5497 13626 5553 13628
rect 5577 13626 5633 13628
rect 5337 13574 5383 13626
rect 5383 13574 5393 13626
rect 5417 13574 5447 13626
rect 5447 13574 5459 13626
rect 5459 13574 5473 13626
rect 5497 13574 5511 13626
rect 5511 13574 5523 13626
rect 5523 13574 5553 13626
rect 5577 13574 5587 13626
rect 5587 13574 5633 13626
rect 5337 13572 5393 13574
rect 5417 13572 5473 13574
rect 5497 13572 5553 13574
rect 5577 13572 5633 13574
rect 3076 13082 3132 13084
rect 3156 13082 3212 13084
rect 3236 13082 3292 13084
rect 3316 13082 3372 13084
rect 3076 13030 3122 13082
rect 3122 13030 3132 13082
rect 3156 13030 3186 13082
rect 3186 13030 3198 13082
rect 3198 13030 3212 13082
rect 3236 13030 3250 13082
rect 3250 13030 3262 13082
rect 3262 13030 3292 13082
rect 3316 13030 3326 13082
rect 3326 13030 3372 13082
rect 3076 13028 3132 13030
rect 3156 13028 3212 13030
rect 3236 13028 3292 13030
rect 3316 13028 3372 13030
rect 2416 12538 2472 12540
rect 2496 12538 2552 12540
rect 2576 12538 2632 12540
rect 2656 12538 2712 12540
rect 2416 12486 2462 12538
rect 2462 12486 2472 12538
rect 2496 12486 2526 12538
rect 2526 12486 2538 12538
rect 2538 12486 2552 12538
rect 2576 12486 2590 12538
rect 2590 12486 2602 12538
rect 2602 12486 2632 12538
rect 2656 12486 2666 12538
rect 2666 12486 2712 12538
rect 2416 12484 2472 12486
rect 2496 12484 2552 12486
rect 2576 12484 2632 12486
rect 2656 12484 2712 12486
rect 5337 12538 5393 12540
rect 5417 12538 5473 12540
rect 5497 12538 5553 12540
rect 5577 12538 5633 12540
rect 5337 12486 5383 12538
rect 5383 12486 5393 12538
rect 5417 12486 5447 12538
rect 5447 12486 5459 12538
rect 5459 12486 5473 12538
rect 5497 12486 5511 12538
rect 5511 12486 5523 12538
rect 5523 12486 5553 12538
rect 5577 12486 5587 12538
rect 5587 12486 5633 12538
rect 5337 12484 5393 12486
rect 5417 12484 5473 12486
rect 5497 12484 5553 12486
rect 5577 12484 5633 12486
rect 3076 11994 3132 11996
rect 3156 11994 3212 11996
rect 3236 11994 3292 11996
rect 3316 11994 3372 11996
rect 3076 11942 3122 11994
rect 3122 11942 3132 11994
rect 3156 11942 3186 11994
rect 3186 11942 3198 11994
rect 3198 11942 3212 11994
rect 3236 11942 3250 11994
rect 3250 11942 3262 11994
rect 3262 11942 3292 11994
rect 3316 11942 3326 11994
rect 3326 11942 3372 11994
rect 3076 11940 3132 11942
rect 3156 11940 3212 11942
rect 3236 11940 3292 11942
rect 3316 11940 3372 11942
rect 2416 11450 2472 11452
rect 2496 11450 2552 11452
rect 2576 11450 2632 11452
rect 2656 11450 2712 11452
rect 2416 11398 2462 11450
rect 2462 11398 2472 11450
rect 2496 11398 2526 11450
rect 2526 11398 2538 11450
rect 2538 11398 2552 11450
rect 2576 11398 2590 11450
rect 2590 11398 2602 11450
rect 2602 11398 2632 11450
rect 2656 11398 2666 11450
rect 2666 11398 2712 11450
rect 2416 11396 2472 11398
rect 2496 11396 2552 11398
rect 2576 11396 2632 11398
rect 2656 11396 2712 11398
rect 5337 11450 5393 11452
rect 5417 11450 5473 11452
rect 5497 11450 5553 11452
rect 5577 11450 5633 11452
rect 5337 11398 5383 11450
rect 5383 11398 5393 11450
rect 5417 11398 5447 11450
rect 5447 11398 5459 11450
rect 5459 11398 5473 11450
rect 5497 11398 5511 11450
rect 5511 11398 5523 11450
rect 5523 11398 5553 11450
rect 5577 11398 5587 11450
rect 5587 11398 5633 11450
rect 5337 11396 5393 11398
rect 5417 11396 5473 11398
rect 5497 11396 5553 11398
rect 5577 11396 5633 11398
rect 3076 10906 3132 10908
rect 3156 10906 3212 10908
rect 3236 10906 3292 10908
rect 3316 10906 3372 10908
rect 3076 10854 3122 10906
rect 3122 10854 3132 10906
rect 3156 10854 3186 10906
rect 3186 10854 3198 10906
rect 3198 10854 3212 10906
rect 3236 10854 3250 10906
rect 3250 10854 3262 10906
rect 3262 10854 3292 10906
rect 3316 10854 3326 10906
rect 3326 10854 3372 10906
rect 3076 10852 3132 10854
rect 3156 10852 3212 10854
rect 3236 10852 3292 10854
rect 3316 10852 3372 10854
rect 2416 10362 2472 10364
rect 2496 10362 2552 10364
rect 2576 10362 2632 10364
rect 2656 10362 2712 10364
rect 2416 10310 2462 10362
rect 2462 10310 2472 10362
rect 2496 10310 2526 10362
rect 2526 10310 2538 10362
rect 2538 10310 2552 10362
rect 2576 10310 2590 10362
rect 2590 10310 2602 10362
rect 2602 10310 2632 10362
rect 2656 10310 2666 10362
rect 2666 10310 2712 10362
rect 2416 10308 2472 10310
rect 2496 10308 2552 10310
rect 2576 10308 2632 10310
rect 2656 10308 2712 10310
rect 3076 9818 3132 9820
rect 3156 9818 3212 9820
rect 3236 9818 3292 9820
rect 3316 9818 3372 9820
rect 3076 9766 3122 9818
rect 3122 9766 3132 9818
rect 3156 9766 3186 9818
rect 3186 9766 3198 9818
rect 3198 9766 3212 9818
rect 3236 9766 3250 9818
rect 3250 9766 3262 9818
rect 3262 9766 3292 9818
rect 3316 9766 3326 9818
rect 3326 9766 3372 9818
rect 3076 9764 3132 9766
rect 3156 9764 3212 9766
rect 3236 9764 3292 9766
rect 3316 9764 3372 9766
rect 2416 9274 2472 9276
rect 2496 9274 2552 9276
rect 2576 9274 2632 9276
rect 2656 9274 2712 9276
rect 2416 9222 2462 9274
rect 2462 9222 2472 9274
rect 2496 9222 2526 9274
rect 2526 9222 2538 9274
rect 2538 9222 2552 9274
rect 2576 9222 2590 9274
rect 2590 9222 2602 9274
rect 2602 9222 2632 9274
rect 2656 9222 2666 9274
rect 2666 9222 2712 9274
rect 2416 9220 2472 9222
rect 2496 9220 2552 9222
rect 2576 9220 2632 9222
rect 2656 9220 2712 9222
rect 5337 10362 5393 10364
rect 5417 10362 5473 10364
rect 5497 10362 5553 10364
rect 5577 10362 5633 10364
rect 5337 10310 5383 10362
rect 5383 10310 5393 10362
rect 5417 10310 5447 10362
rect 5447 10310 5459 10362
rect 5459 10310 5473 10362
rect 5497 10310 5511 10362
rect 5511 10310 5523 10362
rect 5523 10310 5553 10362
rect 5577 10310 5587 10362
rect 5587 10310 5633 10362
rect 5337 10308 5393 10310
rect 5417 10308 5473 10310
rect 5497 10308 5553 10310
rect 5577 10308 5633 10310
rect 3076 8730 3132 8732
rect 3156 8730 3212 8732
rect 3236 8730 3292 8732
rect 3316 8730 3372 8732
rect 3076 8678 3122 8730
rect 3122 8678 3132 8730
rect 3156 8678 3186 8730
rect 3186 8678 3198 8730
rect 3198 8678 3212 8730
rect 3236 8678 3250 8730
rect 3250 8678 3262 8730
rect 3262 8678 3292 8730
rect 3316 8678 3326 8730
rect 3326 8678 3372 8730
rect 3076 8676 3132 8678
rect 3156 8676 3212 8678
rect 3236 8676 3292 8678
rect 3316 8676 3372 8678
rect 5337 9274 5393 9276
rect 5417 9274 5473 9276
rect 5497 9274 5553 9276
rect 5577 9274 5633 9276
rect 5337 9222 5383 9274
rect 5383 9222 5393 9274
rect 5417 9222 5447 9274
rect 5447 9222 5459 9274
rect 5459 9222 5473 9274
rect 5497 9222 5511 9274
rect 5511 9222 5523 9274
rect 5523 9222 5553 9274
rect 5577 9222 5587 9274
rect 5587 9222 5633 9274
rect 5337 9220 5393 9222
rect 5417 9220 5473 9222
rect 5497 9220 5553 9222
rect 5577 9220 5633 9222
rect 2416 8186 2472 8188
rect 2496 8186 2552 8188
rect 2576 8186 2632 8188
rect 2656 8186 2712 8188
rect 2416 8134 2462 8186
rect 2462 8134 2472 8186
rect 2496 8134 2526 8186
rect 2526 8134 2538 8186
rect 2538 8134 2552 8186
rect 2576 8134 2590 8186
rect 2590 8134 2602 8186
rect 2602 8134 2632 8186
rect 2656 8134 2666 8186
rect 2666 8134 2712 8186
rect 2416 8132 2472 8134
rect 2496 8132 2552 8134
rect 2576 8132 2632 8134
rect 2656 8132 2712 8134
rect 3076 7642 3132 7644
rect 3156 7642 3212 7644
rect 3236 7642 3292 7644
rect 3316 7642 3372 7644
rect 3076 7590 3122 7642
rect 3122 7590 3132 7642
rect 3156 7590 3186 7642
rect 3186 7590 3198 7642
rect 3198 7590 3212 7642
rect 3236 7590 3250 7642
rect 3250 7590 3262 7642
rect 3262 7590 3292 7642
rect 3316 7590 3326 7642
rect 3326 7590 3372 7642
rect 3076 7588 3132 7590
rect 3156 7588 3212 7590
rect 3236 7588 3292 7590
rect 3316 7588 3372 7590
rect 2416 7098 2472 7100
rect 2496 7098 2552 7100
rect 2576 7098 2632 7100
rect 2656 7098 2712 7100
rect 2416 7046 2462 7098
rect 2462 7046 2472 7098
rect 2496 7046 2526 7098
rect 2526 7046 2538 7098
rect 2538 7046 2552 7098
rect 2576 7046 2590 7098
rect 2590 7046 2602 7098
rect 2602 7046 2632 7098
rect 2656 7046 2666 7098
rect 2666 7046 2712 7098
rect 2416 7044 2472 7046
rect 2496 7044 2552 7046
rect 2576 7044 2632 7046
rect 2656 7044 2712 7046
rect 3076 6554 3132 6556
rect 3156 6554 3212 6556
rect 3236 6554 3292 6556
rect 3316 6554 3372 6556
rect 3076 6502 3122 6554
rect 3122 6502 3132 6554
rect 3156 6502 3186 6554
rect 3186 6502 3198 6554
rect 3198 6502 3212 6554
rect 3236 6502 3250 6554
rect 3250 6502 3262 6554
rect 3262 6502 3292 6554
rect 3316 6502 3326 6554
rect 3326 6502 3372 6554
rect 3076 6500 3132 6502
rect 3156 6500 3212 6502
rect 3236 6500 3292 6502
rect 3316 6500 3372 6502
rect 2416 6010 2472 6012
rect 2496 6010 2552 6012
rect 2576 6010 2632 6012
rect 2656 6010 2712 6012
rect 2416 5958 2462 6010
rect 2462 5958 2472 6010
rect 2496 5958 2526 6010
rect 2526 5958 2538 6010
rect 2538 5958 2552 6010
rect 2576 5958 2590 6010
rect 2590 5958 2602 6010
rect 2602 5958 2632 6010
rect 2656 5958 2666 6010
rect 2666 5958 2712 6010
rect 2416 5956 2472 5958
rect 2496 5956 2552 5958
rect 2576 5956 2632 5958
rect 2656 5956 2712 5958
rect 1490 4120 1546 4176
rect 1582 3068 1584 3088
rect 1584 3068 1636 3088
rect 1636 3068 1638 3088
rect 1582 3032 1638 3068
rect 3698 6160 3754 6216
rect 3076 5466 3132 5468
rect 3156 5466 3212 5468
rect 3236 5466 3292 5468
rect 3316 5466 3372 5468
rect 3076 5414 3122 5466
rect 3122 5414 3132 5466
rect 3156 5414 3186 5466
rect 3186 5414 3198 5466
rect 3198 5414 3212 5466
rect 3236 5414 3250 5466
rect 3250 5414 3262 5466
rect 3262 5414 3292 5466
rect 3316 5414 3326 5466
rect 3326 5414 3372 5466
rect 3076 5412 3132 5414
rect 3156 5412 3212 5414
rect 3236 5412 3292 5414
rect 3316 5412 3372 5414
rect 2416 4922 2472 4924
rect 2496 4922 2552 4924
rect 2576 4922 2632 4924
rect 2656 4922 2712 4924
rect 2416 4870 2462 4922
rect 2462 4870 2472 4922
rect 2496 4870 2526 4922
rect 2526 4870 2538 4922
rect 2538 4870 2552 4922
rect 2576 4870 2590 4922
rect 2590 4870 2602 4922
rect 2602 4870 2632 4922
rect 2656 4870 2666 4922
rect 2666 4870 2712 4922
rect 2416 4868 2472 4870
rect 2496 4868 2552 4870
rect 2576 4868 2632 4870
rect 2656 4868 2712 4870
rect 3076 4378 3132 4380
rect 3156 4378 3212 4380
rect 3236 4378 3292 4380
rect 3316 4378 3372 4380
rect 3076 4326 3122 4378
rect 3122 4326 3132 4378
rect 3156 4326 3186 4378
rect 3186 4326 3198 4378
rect 3198 4326 3212 4378
rect 3236 4326 3250 4378
rect 3250 4326 3262 4378
rect 3262 4326 3292 4378
rect 3316 4326 3326 4378
rect 3326 4326 3372 4378
rect 3076 4324 3132 4326
rect 3156 4324 3212 4326
rect 3236 4324 3292 4326
rect 3316 4324 3372 4326
rect 5337 8186 5393 8188
rect 5417 8186 5473 8188
rect 5497 8186 5553 8188
rect 5577 8186 5633 8188
rect 5337 8134 5383 8186
rect 5383 8134 5393 8186
rect 5417 8134 5447 8186
rect 5447 8134 5459 8186
rect 5459 8134 5473 8186
rect 5497 8134 5511 8186
rect 5511 8134 5523 8186
rect 5523 8134 5553 8186
rect 5577 8134 5587 8186
rect 5587 8134 5633 8186
rect 5337 8132 5393 8134
rect 5417 8132 5473 8134
rect 5497 8132 5553 8134
rect 5577 8132 5633 8134
rect 4158 5244 4160 5264
rect 4160 5244 4212 5264
rect 4212 5244 4214 5264
rect 4158 5208 4214 5244
rect 3882 5072 3938 5128
rect 2416 3834 2472 3836
rect 2496 3834 2552 3836
rect 2576 3834 2632 3836
rect 2656 3834 2712 3836
rect 2416 3782 2462 3834
rect 2462 3782 2472 3834
rect 2496 3782 2526 3834
rect 2526 3782 2538 3834
rect 2538 3782 2552 3834
rect 2576 3782 2590 3834
rect 2590 3782 2602 3834
rect 2602 3782 2632 3834
rect 2656 3782 2666 3834
rect 2666 3782 2712 3834
rect 2416 3780 2472 3782
rect 2496 3780 2552 3782
rect 2576 3780 2632 3782
rect 2656 3780 2712 3782
rect 3054 4120 3110 4176
rect 3076 3290 3132 3292
rect 3156 3290 3212 3292
rect 3236 3290 3292 3292
rect 3316 3290 3372 3292
rect 3076 3238 3122 3290
rect 3122 3238 3132 3290
rect 3156 3238 3186 3290
rect 3186 3238 3198 3290
rect 3198 3238 3212 3290
rect 3236 3238 3250 3290
rect 3250 3238 3262 3290
rect 3262 3238 3292 3290
rect 3316 3238 3326 3290
rect 3326 3238 3372 3290
rect 3076 3236 3132 3238
rect 3156 3236 3212 3238
rect 3236 3236 3292 3238
rect 3316 3236 3372 3238
rect 2416 2746 2472 2748
rect 2496 2746 2552 2748
rect 2576 2746 2632 2748
rect 2656 2746 2712 2748
rect 2416 2694 2462 2746
rect 2462 2694 2472 2746
rect 2496 2694 2526 2746
rect 2526 2694 2538 2746
rect 2538 2694 2552 2746
rect 2576 2694 2590 2746
rect 2590 2694 2602 2746
rect 2602 2694 2632 2746
rect 2656 2694 2666 2746
rect 2666 2694 2712 2746
rect 2416 2692 2472 2694
rect 2496 2692 2552 2694
rect 2576 2692 2632 2694
rect 2656 2692 2712 2694
rect 4158 2760 4214 2816
rect 3076 2202 3132 2204
rect 3156 2202 3212 2204
rect 3236 2202 3292 2204
rect 3316 2202 3372 2204
rect 3076 2150 3122 2202
rect 3122 2150 3132 2202
rect 3156 2150 3186 2202
rect 3186 2150 3198 2202
rect 3198 2150 3212 2202
rect 3236 2150 3250 2202
rect 3250 2150 3262 2202
rect 3262 2150 3292 2202
rect 3316 2150 3326 2202
rect 3326 2150 3372 2202
rect 3076 2148 3132 2150
rect 3156 2148 3212 2150
rect 3236 2148 3292 2150
rect 3316 2148 3372 2150
rect 5337 7098 5393 7100
rect 5417 7098 5473 7100
rect 5497 7098 5553 7100
rect 5577 7098 5633 7100
rect 5337 7046 5383 7098
rect 5383 7046 5393 7098
rect 5417 7046 5447 7098
rect 5447 7046 5459 7098
rect 5459 7046 5473 7098
rect 5497 7046 5511 7098
rect 5511 7046 5523 7098
rect 5523 7046 5553 7098
rect 5577 7046 5587 7098
rect 5587 7046 5633 7098
rect 5337 7044 5393 7046
rect 5417 7044 5473 7046
rect 5497 7044 5553 7046
rect 5577 7044 5633 7046
rect 8258 13626 8314 13628
rect 8338 13626 8394 13628
rect 8418 13626 8474 13628
rect 8498 13626 8554 13628
rect 8258 13574 8304 13626
rect 8304 13574 8314 13626
rect 8338 13574 8368 13626
rect 8368 13574 8380 13626
rect 8380 13574 8394 13626
rect 8418 13574 8432 13626
rect 8432 13574 8444 13626
rect 8444 13574 8474 13626
rect 8498 13574 8508 13626
rect 8508 13574 8554 13626
rect 8258 13572 8314 13574
rect 8338 13572 8394 13574
rect 8418 13572 8474 13574
rect 8498 13572 8554 13574
rect 11179 13626 11235 13628
rect 11259 13626 11315 13628
rect 11339 13626 11395 13628
rect 11419 13626 11475 13628
rect 11179 13574 11225 13626
rect 11225 13574 11235 13626
rect 11259 13574 11289 13626
rect 11289 13574 11301 13626
rect 11301 13574 11315 13626
rect 11339 13574 11353 13626
rect 11353 13574 11365 13626
rect 11365 13574 11395 13626
rect 11419 13574 11429 13626
rect 11429 13574 11475 13626
rect 11179 13572 11235 13574
rect 11259 13572 11315 13574
rect 11339 13572 11395 13574
rect 11419 13572 11475 13574
rect 5997 13082 6053 13084
rect 6077 13082 6133 13084
rect 6157 13082 6213 13084
rect 6237 13082 6293 13084
rect 5997 13030 6043 13082
rect 6043 13030 6053 13082
rect 6077 13030 6107 13082
rect 6107 13030 6119 13082
rect 6119 13030 6133 13082
rect 6157 13030 6171 13082
rect 6171 13030 6183 13082
rect 6183 13030 6213 13082
rect 6237 13030 6247 13082
rect 6247 13030 6293 13082
rect 5997 13028 6053 13030
rect 6077 13028 6133 13030
rect 6157 13028 6213 13030
rect 6237 13028 6293 13030
rect 5997 11994 6053 11996
rect 6077 11994 6133 11996
rect 6157 11994 6213 11996
rect 6237 11994 6293 11996
rect 5997 11942 6043 11994
rect 6043 11942 6053 11994
rect 6077 11942 6107 11994
rect 6107 11942 6119 11994
rect 6119 11942 6133 11994
rect 6157 11942 6171 11994
rect 6171 11942 6183 11994
rect 6183 11942 6213 11994
rect 6237 11942 6247 11994
rect 6247 11942 6293 11994
rect 5997 11940 6053 11942
rect 6077 11940 6133 11942
rect 6157 11940 6213 11942
rect 6237 11940 6293 11942
rect 8918 13082 8974 13084
rect 8998 13082 9054 13084
rect 9078 13082 9134 13084
rect 9158 13082 9214 13084
rect 8918 13030 8964 13082
rect 8964 13030 8974 13082
rect 8998 13030 9028 13082
rect 9028 13030 9040 13082
rect 9040 13030 9054 13082
rect 9078 13030 9092 13082
rect 9092 13030 9104 13082
rect 9104 13030 9134 13082
rect 9158 13030 9168 13082
rect 9168 13030 9214 13082
rect 8918 13028 8974 13030
rect 8998 13028 9054 13030
rect 9078 13028 9134 13030
rect 9158 13028 9214 13030
rect 11839 13082 11895 13084
rect 11919 13082 11975 13084
rect 11999 13082 12055 13084
rect 12079 13082 12135 13084
rect 11839 13030 11885 13082
rect 11885 13030 11895 13082
rect 11919 13030 11949 13082
rect 11949 13030 11961 13082
rect 11961 13030 11975 13082
rect 11999 13030 12013 13082
rect 12013 13030 12025 13082
rect 12025 13030 12055 13082
rect 12079 13030 12089 13082
rect 12089 13030 12135 13082
rect 11839 13028 11895 13030
rect 11919 13028 11975 13030
rect 11999 13028 12055 13030
rect 12079 13028 12135 13030
rect 5997 10906 6053 10908
rect 6077 10906 6133 10908
rect 6157 10906 6213 10908
rect 6237 10906 6293 10908
rect 5997 10854 6043 10906
rect 6043 10854 6053 10906
rect 6077 10854 6107 10906
rect 6107 10854 6119 10906
rect 6119 10854 6133 10906
rect 6157 10854 6171 10906
rect 6171 10854 6183 10906
rect 6183 10854 6213 10906
rect 6237 10854 6247 10906
rect 6247 10854 6293 10906
rect 5997 10852 6053 10854
rect 6077 10852 6133 10854
rect 6157 10852 6213 10854
rect 6237 10852 6293 10854
rect 8258 12538 8314 12540
rect 8338 12538 8394 12540
rect 8418 12538 8474 12540
rect 8498 12538 8554 12540
rect 8258 12486 8304 12538
rect 8304 12486 8314 12538
rect 8338 12486 8368 12538
rect 8368 12486 8380 12538
rect 8380 12486 8394 12538
rect 8418 12486 8432 12538
rect 8432 12486 8444 12538
rect 8444 12486 8474 12538
rect 8498 12486 8508 12538
rect 8508 12486 8554 12538
rect 8258 12484 8314 12486
rect 8338 12484 8394 12486
rect 8418 12484 8474 12486
rect 8498 12484 8554 12486
rect 11179 12538 11235 12540
rect 11259 12538 11315 12540
rect 11339 12538 11395 12540
rect 11419 12538 11475 12540
rect 11179 12486 11225 12538
rect 11225 12486 11235 12538
rect 11259 12486 11289 12538
rect 11289 12486 11301 12538
rect 11301 12486 11315 12538
rect 11339 12486 11353 12538
rect 11353 12486 11365 12538
rect 11365 12486 11395 12538
rect 11419 12486 11429 12538
rect 11429 12486 11475 12538
rect 11179 12484 11235 12486
rect 11259 12484 11315 12486
rect 11339 12484 11395 12486
rect 11419 12484 11475 12486
rect 8918 11994 8974 11996
rect 8998 11994 9054 11996
rect 9078 11994 9134 11996
rect 9158 11994 9214 11996
rect 8918 11942 8964 11994
rect 8964 11942 8974 11994
rect 8998 11942 9028 11994
rect 9028 11942 9040 11994
rect 9040 11942 9054 11994
rect 9078 11942 9092 11994
rect 9092 11942 9104 11994
rect 9104 11942 9134 11994
rect 9158 11942 9168 11994
rect 9168 11942 9214 11994
rect 8918 11940 8974 11942
rect 8998 11940 9054 11942
rect 9078 11940 9134 11942
rect 9158 11940 9214 11942
rect 11839 11994 11895 11996
rect 11919 11994 11975 11996
rect 11999 11994 12055 11996
rect 12079 11994 12135 11996
rect 11839 11942 11885 11994
rect 11885 11942 11895 11994
rect 11919 11942 11949 11994
rect 11949 11942 11961 11994
rect 11961 11942 11975 11994
rect 11999 11942 12013 11994
rect 12013 11942 12025 11994
rect 12025 11942 12055 11994
rect 12079 11942 12089 11994
rect 12089 11942 12135 11994
rect 11839 11940 11895 11942
rect 11919 11940 11975 11942
rect 11999 11940 12055 11942
rect 12079 11940 12135 11942
rect 8258 11450 8314 11452
rect 8338 11450 8394 11452
rect 8418 11450 8474 11452
rect 8498 11450 8554 11452
rect 8258 11398 8304 11450
rect 8304 11398 8314 11450
rect 8338 11398 8368 11450
rect 8368 11398 8380 11450
rect 8380 11398 8394 11450
rect 8418 11398 8432 11450
rect 8432 11398 8444 11450
rect 8444 11398 8474 11450
rect 8498 11398 8508 11450
rect 8508 11398 8554 11450
rect 8258 11396 8314 11398
rect 8338 11396 8394 11398
rect 8418 11396 8474 11398
rect 8498 11396 8554 11398
rect 11179 11450 11235 11452
rect 11259 11450 11315 11452
rect 11339 11450 11395 11452
rect 11419 11450 11475 11452
rect 11179 11398 11225 11450
rect 11225 11398 11235 11450
rect 11259 11398 11289 11450
rect 11289 11398 11301 11450
rect 11301 11398 11315 11450
rect 11339 11398 11353 11450
rect 11353 11398 11365 11450
rect 11365 11398 11395 11450
rect 11419 11398 11429 11450
rect 11429 11398 11475 11450
rect 11179 11396 11235 11398
rect 11259 11396 11315 11398
rect 11339 11396 11395 11398
rect 11419 11396 11475 11398
rect 8918 10906 8974 10908
rect 8998 10906 9054 10908
rect 9078 10906 9134 10908
rect 9158 10906 9214 10908
rect 8918 10854 8964 10906
rect 8964 10854 8974 10906
rect 8998 10854 9028 10906
rect 9028 10854 9040 10906
rect 9040 10854 9054 10906
rect 9078 10854 9092 10906
rect 9092 10854 9104 10906
rect 9104 10854 9134 10906
rect 9158 10854 9168 10906
rect 9168 10854 9214 10906
rect 8918 10852 8974 10854
rect 8998 10852 9054 10854
rect 9078 10852 9134 10854
rect 9158 10852 9214 10854
rect 11839 10906 11895 10908
rect 11919 10906 11975 10908
rect 11999 10906 12055 10908
rect 12079 10906 12135 10908
rect 11839 10854 11885 10906
rect 11885 10854 11895 10906
rect 11919 10854 11949 10906
rect 11949 10854 11961 10906
rect 11961 10854 11975 10906
rect 11999 10854 12013 10906
rect 12013 10854 12025 10906
rect 12025 10854 12055 10906
rect 12079 10854 12089 10906
rect 12089 10854 12135 10906
rect 11839 10852 11895 10854
rect 11919 10852 11975 10854
rect 11999 10852 12055 10854
rect 12079 10852 12135 10854
rect 8258 10362 8314 10364
rect 8338 10362 8394 10364
rect 8418 10362 8474 10364
rect 8498 10362 8554 10364
rect 8258 10310 8304 10362
rect 8304 10310 8314 10362
rect 8338 10310 8368 10362
rect 8368 10310 8380 10362
rect 8380 10310 8394 10362
rect 8418 10310 8432 10362
rect 8432 10310 8444 10362
rect 8444 10310 8474 10362
rect 8498 10310 8508 10362
rect 8508 10310 8554 10362
rect 8258 10308 8314 10310
rect 8338 10308 8394 10310
rect 8418 10308 8474 10310
rect 8498 10308 8554 10310
rect 11179 10362 11235 10364
rect 11259 10362 11315 10364
rect 11339 10362 11395 10364
rect 11419 10362 11475 10364
rect 11179 10310 11225 10362
rect 11225 10310 11235 10362
rect 11259 10310 11289 10362
rect 11289 10310 11301 10362
rect 11301 10310 11315 10362
rect 11339 10310 11353 10362
rect 11353 10310 11365 10362
rect 11365 10310 11395 10362
rect 11419 10310 11429 10362
rect 11429 10310 11475 10362
rect 11179 10308 11235 10310
rect 11259 10308 11315 10310
rect 11339 10308 11395 10310
rect 11419 10308 11475 10310
rect 5997 9818 6053 9820
rect 6077 9818 6133 9820
rect 6157 9818 6213 9820
rect 6237 9818 6293 9820
rect 5997 9766 6043 9818
rect 6043 9766 6053 9818
rect 6077 9766 6107 9818
rect 6107 9766 6119 9818
rect 6119 9766 6133 9818
rect 6157 9766 6171 9818
rect 6171 9766 6183 9818
rect 6183 9766 6213 9818
rect 6237 9766 6247 9818
rect 6247 9766 6293 9818
rect 5997 9764 6053 9766
rect 6077 9764 6133 9766
rect 6157 9764 6213 9766
rect 6237 9764 6293 9766
rect 5997 8730 6053 8732
rect 6077 8730 6133 8732
rect 6157 8730 6213 8732
rect 6237 8730 6293 8732
rect 5997 8678 6043 8730
rect 6043 8678 6053 8730
rect 6077 8678 6107 8730
rect 6107 8678 6119 8730
rect 6119 8678 6133 8730
rect 6157 8678 6171 8730
rect 6171 8678 6183 8730
rect 6183 8678 6213 8730
rect 6237 8678 6247 8730
rect 6247 8678 6293 8730
rect 5997 8676 6053 8678
rect 6077 8676 6133 8678
rect 6157 8676 6213 8678
rect 6237 8676 6293 8678
rect 5997 7642 6053 7644
rect 6077 7642 6133 7644
rect 6157 7642 6213 7644
rect 6237 7642 6293 7644
rect 5997 7590 6043 7642
rect 6043 7590 6053 7642
rect 6077 7590 6107 7642
rect 6107 7590 6119 7642
rect 6119 7590 6133 7642
rect 6157 7590 6171 7642
rect 6171 7590 6183 7642
rect 6183 7590 6213 7642
rect 6237 7590 6247 7642
rect 6247 7590 6293 7642
rect 5997 7588 6053 7590
rect 6077 7588 6133 7590
rect 6157 7588 6213 7590
rect 6237 7588 6293 7590
rect 5337 6010 5393 6012
rect 5417 6010 5473 6012
rect 5497 6010 5553 6012
rect 5577 6010 5633 6012
rect 5337 5958 5383 6010
rect 5383 5958 5393 6010
rect 5417 5958 5447 6010
rect 5447 5958 5459 6010
rect 5459 5958 5473 6010
rect 5497 5958 5511 6010
rect 5511 5958 5523 6010
rect 5523 5958 5553 6010
rect 5577 5958 5587 6010
rect 5587 5958 5633 6010
rect 5337 5956 5393 5958
rect 5417 5956 5473 5958
rect 5497 5956 5553 5958
rect 5577 5956 5633 5958
rect 5078 4140 5134 4176
rect 5078 4120 5080 4140
rect 5080 4120 5132 4140
rect 5132 4120 5134 4140
rect 4710 3476 4712 3496
rect 4712 3476 4764 3496
rect 4764 3476 4766 3496
rect 4710 3440 4766 3476
rect 4434 3052 4490 3088
rect 4434 3032 4436 3052
rect 4436 3032 4488 3052
rect 4488 3032 4490 3052
rect 4986 3576 5042 3632
rect 5337 4922 5393 4924
rect 5417 4922 5473 4924
rect 5497 4922 5553 4924
rect 5577 4922 5633 4924
rect 5337 4870 5383 4922
rect 5383 4870 5393 4922
rect 5417 4870 5447 4922
rect 5447 4870 5459 4922
rect 5459 4870 5473 4922
rect 5497 4870 5511 4922
rect 5511 4870 5523 4922
rect 5523 4870 5553 4922
rect 5577 4870 5587 4922
rect 5587 4870 5633 4922
rect 5337 4868 5393 4870
rect 5417 4868 5473 4870
rect 5497 4868 5553 4870
rect 5577 4868 5633 4870
rect 5997 6554 6053 6556
rect 6077 6554 6133 6556
rect 6157 6554 6213 6556
rect 6237 6554 6293 6556
rect 5997 6502 6043 6554
rect 6043 6502 6053 6554
rect 6077 6502 6107 6554
rect 6107 6502 6119 6554
rect 6119 6502 6133 6554
rect 6157 6502 6171 6554
rect 6171 6502 6183 6554
rect 6183 6502 6213 6554
rect 6237 6502 6247 6554
rect 6247 6502 6293 6554
rect 5997 6500 6053 6502
rect 6077 6500 6133 6502
rect 6157 6500 6213 6502
rect 6237 6500 6293 6502
rect 6182 6160 6238 6216
rect 5997 5466 6053 5468
rect 6077 5466 6133 5468
rect 6157 5466 6213 5468
rect 6237 5466 6293 5468
rect 5997 5414 6043 5466
rect 6043 5414 6053 5466
rect 6077 5414 6107 5466
rect 6107 5414 6119 5466
rect 6119 5414 6133 5466
rect 6157 5414 6171 5466
rect 6171 5414 6183 5466
rect 6183 5414 6213 5466
rect 6237 5414 6247 5466
rect 6247 5414 6293 5466
rect 5997 5412 6053 5414
rect 6077 5412 6133 5414
rect 6157 5412 6213 5414
rect 6237 5412 6293 5414
rect 6274 5228 6330 5264
rect 6274 5208 6276 5228
rect 6276 5208 6328 5228
rect 6328 5208 6330 5228
rect 5997 4378 6053 4380
rect 6077 4378 6133 4380
rect 6157 4378 6213 4380
rect 6237 4378 6293 4380
rect 5997 4326 6043 4378
rect 6043 4326 6053 4378
rect 6077 4326 6107 4378
rect 6107 4326 6119 4378
rect 6119 4326 6133 4378
rect 6157 4326 6171 4378
rect 6171 4326 6183 4378
rect 6183 4326 6213 4378
rect 6237 4326 6247 4378
rect 6247 4326 6293 4378
rect 5997 4324 6053 4326
rect 6077 4324 6133 4326
rect 6157 4324 6213 4326
rect 6237 4324 6293 4326
rect 5722 4120 5778 4176
rect 5337 3834 5393 3836
rect 5417 3834 5473 3836
rect 5497 3834 5553 3836
rect 5577 3834 5633 3836
rect 5337 3782 5383 3834
rect 5383 3782 5393 3834
rect 5417 3782 5447 3834
rect 5447 3782 5459 3834
rect 5459 3782 5473 3834
rect 5497 3782 5511 3834
rect 5511 3782 5523 3834
rect 5523 3782 5553 3834
rect 5577 3782 5587 3834
rect 5587 3782 5633 3834
rect 5337 3780 5393 3782
rect 5417 3780 5473 3782
rect 5497 3780 5553 3782
rect 5577 3780 5633 3782
rect 4894 2896 4950 2952
rect 5078 2760 5134 2816
rect 5337 2746 5393 2748
rect 5417 2746 5473 2748
rect 5497 2746 5553 2748
rect 5577 2746 5633 2748
rect 5337 2694 5383 2746
rect 5383 2694 5393 2746
rect 5417 2694 5447 2746
rect 5447 2694 5459 2746
rect 5459 2694 5473 2746
rect 5497 2694 5511 2746
rect 5511 2694 5523 2746
rect 5523 2694 5553 2746
rect 5577 2694 5587 2746
rect 5587 2694 5633 2746
rect 5337 2692 5393 2694
rect 5417 2692 5473 2694
rect 5497 2692 5553 2694
rect 5577 2692 5633 2694
rect 5997 3290 6053 3292
rect 6077 3290 6133 3292
rect 6157 3290 6213 3292
rect 6237 3290 6293 3292
rect 5997 3238 6043 3290
rect 6043 3238 6053 3290
rect 6077 3238 6107 3290
rect 6107 3238 6119 3290
rect 6119 3238 6133 3290
rect 6157 3238 6171 3290
rect 6171 3238 6183 3290
rect 6183 3238 6213 3290
rect 6237 3238 6247 3290
rect 6247 3238 6293 3290
rect 5997 3236 6053 3238
rect 6077 3236 6133 3238
rect 6157 3236 6213 3238
rect 6237 3236 6293 3238
rect 7562 6160 7618 6216
rect 6918 5228 6974 5264
rect 6918 5208 6920 5228
rect 6920 5208 6972 5228
rect 6972 5208 6974 5228
rect 7102 5092 7158 5128
rect 7102 5072 7104 5092
rect 7104 5072 7156 5092
rect 7156 5072 7158 5092
rect 8918 9818 8974 9820
rect 8998 9818 9054 9820
rect 9078 9818 9134 9820
rect 9158 9818 9214 9820
rect 8918 9766 8964 9818
rect 8964 9766 8974 9818
rect 8998 9766 9028 9818
rect 9028 9766 9040 9818
rect 9040 9766 9054 9818
rect 9078 9766 9092 9818
rect 9092 9766 9104 9818
rect 9104 9766 9134 9818
rect 9158 9766 9168 9818
rect 9168 9766 9214 9818
rect 8918 9764 8974 9766
rect 8998 9764 9054 9766
rect 9078 9764 9134 9766
rect 9158 9764 9214 9766
rect 11839 9818 11895 9820
rect 11919 9818 11975 9820
rect 11999 9818 12055 9820
rect 12079 9818 12135 9820
rect 11839 9766 11885 9818
rect 11885 9766 11895 9818
rect 11919 9766 11949 9818
rect 11949 9766 11961 9818
rect 11961 9766 11975 9818
rect 11999 9766 12013 9818
rect 12013 9766 12025 9818
rect 12025 9766 12055 9818
rect 12079 9766 12089 9818
rect 12089 9766 12135 9818
rect 11839 9764 11895 9766
rect 11919 9764 11975 9766
rect 11999 9764 12055 9766
rect 12079 9764 12135 9766
rect 8258 9274 8314 9276
rect 8338 9274 8394 9276
rect 8418 9274 8474 9276
rect 8498 9274 8554 9276
rect 8258 9222 8304 9274
rect 8304 9222 8314 9274
rect 8338 9222 8368 9274
rect 8368 9222 8380 9274
rect 8380 9222 8394 9274
rect 8418 9222 8432 9274
rect 8432 9222 8444 9274
rect 8444 9222 8474 9274
rect 8498 9222 8508 9274
rect 8508 9222 8554 9274
rect 8258 9220 8314 9222
rect 8338 9220 8394 9222
rect 8418 9220 8474 9222
rect 8498 9220 8554 9222
rect 11179 9274 11235 9276
rect 11259 9274 11315 9276
rect 11339 9274 11395 9276
rect 11419 9274 11475 9276
rect 11179 9222 11225 9274
rect 11225 9222 11235 9274
rect 11259 9222 11289 9274
rect 11289 9222 11301 9274
rect 11301 9222 11315 9274
rect 11339 9222 11353 9274
rect 11353 9222 11365 9274
rect 11365 9222 11395 9274
rect 11419 9222 11429 9274
rect 11429 9222 11475 9274
rect 11179 9220 11235 9222
rect 11259 9220 11315 9222
rect 11339 9220 11395 9222
rect 11419 9220 11475 9222
rect 8918 8730 8974 8732
rect 8998 8730 9054 8732
rect 9078 8730 9134 8732
rect 9158 8730 9214 8732
rect 8918 8678 8964 8730
rect 8964 8678 8974 8730
rect 8998 8678 9028 8730
rect 9028 8678 9040 8730
rect 9040 8678 9054 8730
rect 9078 8678 9092 8730
rect 9092 8678 9104 8730
rect 9104 8678 9134 8730
rect 9158 8678 9168 8730
rect 9168 8678 9214 8730
rect 8918 8676 8974 8678
rect 8998 8676 9054 8678
rect 9078 8676 9134 8678
rect 9158 8676 9214 8678
rect 8258 8186 8314 8188
rect 8338 8186 8394 8188
rect 8418 8186 8474 8188
rect 8498 8186 8554 8188
rect 8258 8134 8304 8186
rect 8304 8134 8314 8186
rect 8338 8134 8368 8186
rect 8368 8134 8380 8186
rect 8380 8134 8394 8186
rect 8418 8134 8432 8186
rect 8432 8134 8444 8186
rect 8444 8134 8474 8186
rect 8498 8134 8508 8186
rect 8508 8134 8554 8186
rect 8258 8132 8314 8134
rect 8338 8132 8394 8134
rect 8418 8132 8474 8134
rect 8498 8132 8554 8134
rect 11839 8730 11895 8732
rect 11919 8730 11975 8732
rect 11999 8730 12055 8732
rect 12079 8730 12135 8732
rect 11839 8678 11885 8730
rect 11885 8678 11895 8730
rect 11919 8678 11949 8730
rect 11949 8678 11961 8730
rect 11961 8678 11975 8730
rect 11999 8678 12013 8730
rect 12013 8678 12025 8730
rect 12025 8678 12055 8730
rect 12079 8678 12089 8730
rect 12089 8678 12135 8730
rect 11839 8676 11895 8678
rect 11919 8676 11975 8678
rect 11999 8676 12055 8678
rect 12079 8676 12135 8678
rect 11179 8186 11235 8188
rect 11259 8186 11315 8188
rect 11339 8186 11395 8188
rect 11419 8186 11475 8188
rect 11179 8134 11225 8186
rect 11225 8134 11235 8186
rect 11259 8134 11289 8186
rect 11289 8134 11301 8186
rect 11301 8134 11315 8186
rect 11339 8134 11353 8186
rect 11353 8134 11365 8186
rect 11365 8134 11395 8186
rect 11419 8134 11429 8186
rect 11429 8134 11475 8186
rect 11179 8132 11235 8134
rect 11259 8132 11315 8134
rect 11339 8132 11395 8134
rect 11419 8132 11475 8134
rect 8918 7642 8974 7644
rect 8998 7642 9054 7644
rect 9078 7642 9134 7644
rect 9158 7642 9214 7644
rect 8918 7590 8964 7642
rect 8964 7590 8974 7642
rect 8998 7590 9028 7642
rect 9028 7590 9040 7642
rect 9040 7590 9054 7642
rect 9078 7590 9092 7642
rect 9092 7590 9104 7642
rect 9104 7590 9134 7642
rect 9158 7590 9168 7642
rect 9168 7590 9214 7642
rect 8918 7588 8974 7590
rect 8998 7588 9054 7590
rect 9078 7588 9134 7590
rect 9158 7588 9214 7590
rect 11839 7642 11895 7644
rect 11919 7642 11975 7644
rect 11999 7642 12055 7644
rect 12079 7642 12135 7644
rect 11839 7590 11885 7642
rect 11885 7590 11895 7642
rect 11919 7590 11949 7642
rect 11949 7590 11961 7642
rect 11961 7590 11975 7642
rect 11999 7590 12013 7642
rect 12013 7590 12025 7642
rect 12025 7590 12055 7642
rect 12079 7590 12089 7642
rect 12089 7590 12135 7642
rect 11839 7588 11895 7590
rect 11919 7588 11975 7590
rect 11999 7588 12055 7590
rect 12079 7588 12135 7590
rect 8258 7098 8314 7100
rect 8338 7098 8394 7100
rect 8418 7098 8474 7100
rect 8498 7098 8554 7100
rect 8258 7046 8304 7098
rect 8304 7046 8314 7098
rect 8338 7046 8368 7098
rect 8368 7046 8380 7098
rect 8380 7046 8394 7098
rect 8418 7046 8432 7098
rect 8432 7046 8444 7098
rect 8444 7046 8474 7098
rect 8498 7046 8508 7098
rect 8508 7046 8554 7098
rect 8258 7044 8314 7046
rect 8338 7044 8394 7046
rect 8418 7044 8474 7046
rect 8498 7044 8554 7046
rect 7746 5652 7748 5672
rect 7748 5652 7800 5672
rect 7800 5652 7802 5672
rect 7746 5616 7802 5652
rect 8574 6296 8630 6352
rect 7010 3576 7066 3632
rect 8258 6010 8314 6012
rect 8338 6010 8394 6012
rect 8418 6010 8474 6012
rect 8498 6010 8554 6012
rect 8258 5958 8304 6010
rect 8304 5958 8314 6010
rect 8338 5958 8368 6010
rect 8368 5958 8380 6010
rect 8380 5958 8394 6010
rect 8418 5958 8432 6010
rect 8432 5958 8444 6010
rect 8444 5958 8474 6010
rect 8498 5958 8508 6010
rect 8508 5958 8554 6010
rect 8258 5956 8314 5958
rect 8338 5956 8394 5958
rect 8418 5956 8474 5958
rect 8498 5956 8554 5958
rect 8918 6554 8974 6556
rect 8998 6554 9054 6556
rect 9078 6554 9134 6556
rect 9158 6554 9214 6556
rect 8918 6502 8964 6554
rect 8964 6502 8974 6554
rect 8998 6502 9028 6554
rect 9028 6502 9040 6554
rect 9040 6502 9054 6554
rect 9078 6502 9092 6554
rect 9092 6502 9104 6554
rect 9104 6502 9134 6554
rect 9158 6502 9168 6554
rect 9168 6502 9214 6554
rect 8918 6500 8974 6502
rect 8998 6500 9054 6502
rect 9078 6500 9134 6502
rect 9158 6500 9214 6502
rect 9034 6316 9090 6352
rect 9034 6296 9036 6316
rect 9036 6296 9088 6316
rect 9088 6296 9090 6316
rect 8942 6160 8998 6216
rect 8390 5072 8446 5128
rect 8258 4922 8314 4924
rect 8338 4922 8394 4924
rect 8418 4922 8474 4924
rect 8498 4922 8554 4924
rect 8258 4870 8304 4922
rect 8304 4870 8314 4922
rect 8338 4870 8368 4922
rect 8368 4870 8380 4922
rect 8380 4870 8394 4922
rect 8418 4870 8432 4922
rect 8432 4870 8444 4922
rect 8444 4870 8474 4922
rect 8498 4870 8508 4922
rect 8508 4870 8554 4922
rect 8258 4868 8314 4870
rect 8338 4868 8394 4870
rect 8418 4868 8474 4870
rect 8498 4868 8554 4870
rect 7930 4156 7932 4176
rect 7932 4156 7984 4176
rect 7984 4156 7986 4176
rect 7930 4120 7986 4156
rect 8258 3834 8314 3836
rect 8338 3834 8394 3836
rect 8418 3834 8474 3836
rect 8498 3834 8554 3836
rect 8258 3782 8304 3834
rect 8304 3782 8314 3834
rect 8338 3782 8368 3834
rect 8368 3782 8380 3834
rect 8380 3782 8394 3834
rect 8418 3782 8432 3834
rect 8432 3782 8444 3834
rect 8444 3782 8474 3834
rect 8498 3782 8508 3834
rect 8508 3782 8554 3834
rect 8258 3780 8314 3782
rect 8338 3780 8394 3782
rect 8418 3780 8474 3782
rect 8498 3780 8554 3782
rect 9310 5616 9366 5672
rect 8918 5466 8974 5468
rect 8998 5466 9054 5468
rect 9078 5466 9134 5468
rect 9158 5466 9214 5468
rect 8918 5414 8964 5466
rect 8964 5414 8974 5466
rect 8998 5414 9028 5466
rect 9028 5414 9040 5466
rect 9040 5414 9054 5466
rect 9078 5414 9092 5466
rect 9092 5414 9104 5466
rect 9104 5414 9134 5466
rect 9158 5414 9168 5466
rect 9168 5414 9214 5466
rect 8918 5412 8974 5414
rect 8998 5412 9054 5414
rect 9078 5412 9134 5414
rect 9158 5412 9214 5414
rect 8942 4528 8998 4584
rect 8918 4378 8974 4380
rect 8998 4378 9054 4380
rect 9078 4378 9134 4380
rect 9158 4378 9214 4380
rect 8918 4326 8964 4378
rect 8964 4326 8974 4378
rect 8998 4326 9028 4378
rect 9028 4326 9040 4378
rect 9040 4326 9054 4378
rect 9078 4326 9092 4378
rect 9092 4326 9104 4378
rect 9104 4326 9134 4378
rect 9158 4326 9168 4378
rect 9168 4326 9214 4378
rect 8918 4324 8974 4326
rect 8998 4324 9054 4326
rect 9078 4324 9134 4326
rect 9158 4324 9214 4326
rect 7930 3476 7932 3496
rect 7932 3476 7984 3496
rect 7984 3476 7986 3496
rect 7930 3440 7986 3476
rect 8258 2746 8314 2748
rect 8338 2746 8394 2748
rect 8418 2746 8474 2748
rect 8498 2746 8554 2748
rect 8258 2694 8304 2746
rect 8304 2694 8314 2746
rect 8338 2694 8368 2746
rect 8368 2694 8380 2746
rect 8380 2694 8394 2746
rect 8418 2694 8432 2746
rect 8432 2694 8444 2746
rect 8444 2694 8474 2746
rect 8498 2694 8508 2746
rect 8508 2694 8554 2746
rect 8258 2692 8314 2694
rect 8338 2692 8394 2694
rect 8418 2692 8474 2694
rect 8498 2692 8554 2694
rect 9678 6160 9734 6216
rect 11179 7098 11235 7100
rect 11259 7098 11315 7100
rect 11339 7098 11395 7100
rect 11419 7098 11475 7100
rect 11179 7046 11225 7098
rect 11225 7046 11235 7098
rect 11259 7046 11289 7098
rect 11289 7046 11301 7098
rect 11301 7046 11315 7098
rect 11339 7046 11353 7098
rect 11353 7046 11365 7098
rect 11365 7046 11395 7098
rect 11419 7046 11429 7098
rect 11429 7046 11475 7098
rect 11179 7044 11235 7046
rect 11259 7044 11315 7046
rect 11339 7044 11395 7046
rect 11419 7044 11475 7046
rect 11839 6554 11895 6556
rect 11919 6554 11975 6556
rect 11999 6554 12055 6556
rect 12079 6554 12135 6556
rect 11839 6502 11885 6554
rect 11885 6502 11895 6554
rect 11919 6502 11949 6554
rect 11949 6502 11961 6554
rect 11961 6502 11975 6554
rect 11999 6502 12013 6554
rect 12013 6502 12025 6554
rect 12025 6502 12055 6554
rect 12079 6502 12089 6554
rect 12089 6502 12135 6554
rect 11839 6500 11895 6502
rect 11919 6500 11975 6502
rect 11999 6500 12055 6502
rect 12079 6500 12135 6502
rect 9402 4256 9458 4312
rect 8918 3290 8974 3292
rect 8998 3290 9054 3292
rect 9078 3290 9134 3292
rect 9158 3290 9214 3292
rect 8918 3238 8964 3290
rect 8964 3238 8974 3290
rect 8998 3238 9028 3290
rect 9028 3238 9040 3290
rect 9040 3238 9054 3290
rect 9078 3238 9092 3290
rect 9092 3238 9104 3290
rect 9104 3238 9134 3290
rect 9158 3238 9168 3290
rect 9168 3238 9214 3290
rect 8918 3236 8974 3238
rect 8998 3236 9054 3238
rect 9078 3236 9134 3238
rect 9158 3236 9214 3238
rect 9034 2896 9090 2952
rect 10230 6196 10232 6216
rect 10232 6196 10284 6216
rect 10284 6196 10286 6216
rect 10230 6160 10286 6196
rect 11179 6010 11235 6012
rect 11259 6010 11315 6012
rect 11339 6010 11395 6012
rect 11419 6010 11475 6012
rect 11179 5958 11225 6010
rect 11225 5958 11235 6010
rect 11259 5958 11289 6010
rect 11289 5958 11301 6010
rect 11301 5958 11315 6010
rect 11339 5958 11353 6010
rect 11353 5958 11365 6010
rect 11365 5958 11395 6010
rect 11419 5958 11429 6010
rect 11429 5958 11475 6010
rect 11179 5956 11235 5958
rect 11259 5956 11315 5958
rect 11339 5956 11395 5958
rect 11419 5956 11475 5958
rect 11839 5466 11895 5468
rect 11919 5466 11975 5468
rect 11999 5466 12055 5468
rect 12079 5466 12135 5468
rect 11839 5414 11885 5466
rect 11885 5414 11895 5466
rect 11919 5414 11949 5466
rect 11949 5414 11961 5466
rect 11961 5414 11975 5466
rect 11999 5414 12013 5466
rect 12013 5414 12025 5466
rect 12025 5414 12055 5466
rect 12079 5414 12089 5466
rect 12089 5414 12135 5466
rect 11839 5412 11895 5414
rect 11919 5412 11975 5414
rect 11999 5412 12055 5414
rect 12079 5412 12135 5414
rect 11179 4922 11235 4924
rect 11259 4922 11315 4924
rect 11339 4922 11395 4924
rect 11419 4922 11475 4924
rect 11179 4870 11225 4922
rect 11225 4870 11235 4922
rect 11259 4870 11289 4922
rect 11289 4870 11301 4922
rect 11301 4870 11315 4922
rect 11339 4870 11353 4922
rect 11353 4870 11365 4922
rect 11365 4870 11395 4922
rect 11419 4870 11429 4922
rect 11429 4870 11475 4922
rect 11179 4868 11235 4870
rect 11259 4868 11315 4870
rect 11339 4868 11395 4870
rect 11419 4868 11475 4870
rect 11839 4378 11895 4380
rect 11919 4378 11975 4380
rect 11999 4378 12055 4380
rect 12079 4378 12135 4380
rect 11839 4326 11885 4378
rect 11885 4326 11895 4378
rect 11919 4326 11949 4378
rect 11949 4326 11961 4378
rect 11961 4326 11975 4378
rect 11999 4326 12013 4378
rect 12013 4326 12025 4378
rect 12025 4326 12055 4378
rect 12079 4326 12089 4378
rect 12089 4326 12135 4378
rect 11839 4324 11895 4326
rect 11919 4324 11975 4326
rect 11999 4324 12055 4326
rect 12079 4324 12135 4326
rect 11179 3834 11235 3836
rect 11259 3834 11315 3836
rect 11339 3834 11395 3836
rect 11419 3834 11475 3836
rect 11179 3782 11225 3834
rect 11225 3782 11235 3834
rect 11259 3782 11289 3834
rect 11289 3782 11301 3834
rect 11301 3782 11315 3834
rect 11339 3782 11353 3834
rect 11353 3782 11365 3834
rect 11365 3782 11395 3834
rect 11419 3782 11429 3834
rect 11429 3782 11475 3834
rect 11179 3780 11235 3782
rect 11259 3780 11315 3782
rect 11339 3780 11395 3782
rect 11419 3780 11475 3782
rect 11839 3290 11895 3292
rect 11919 3290 11975 3292
rect 11999 3290 12055 3292
rect 12079 3290 12135 3292
rect 11839 3238 11885 3290
rect 11885 3238 11895 3290
rect 11919 3238 11949 3290
rect 11949 3238 11961 3290
rect 11961 3238 11975 3290
rect 11999 3238 12013 3290
rect 12013 3238 12025 3290
rect 12025 3238 12055 3290
rect 12079 3238 12089 3290
rect 12089 3238 12135 3290
rect 11839 3236 11895 3238
rect 11919 3236 11975 3238
rect 11999 3236 12055 3238
rect 12079 3236 12135 3238
rect 11179 2746 11235 2748
rect 11259 2746 11315 2748
rect 11339 2746 11395 2748
rect 11419 2746 11475 2748
rect 11179 2694 11225 2746
rect 11225 2694 11235 2746
rect 11259 2694 11289 2746
rect 11289 2694 11301 2746
rect 11301 2694 11315 2746
rect 11339 2694 11353 2746
rect 11353 2694 11365 2746
rect 11365 2694 11395 2746
rect 11419 2694 11429 2746
rect 11429 2694 11475 2746
rect 11179 2692 11235 2694
rect 11259 2692 11315 2694
rect 11339 2692 11395 2694
rect 11419 2692 11475 2694
rect 5997 2202 6053 2204
rect 6077 2202 6133 2204
rect 6157 2202 6213 2204
rect 6237 2202 6293 2204
rect 5997 2150 6043 2202
rect 6043 2150 6053 2202
rect 6077 2150 6107 2202
rect 6107 2150 6119 2202
rect 6119 2150 6133 2202
rect 6157 2150 6171 2202
rect 6171 2150 6183 2202
rect 6183 2150 6213 2202
rect 6237 2150 6247 2202
rect 6247 2150 6293 2202
rect 5997 2148 6053 2150
rect 6077 2148 6133 2150
rect 6157 2148 6213 2150
rect 6237 2148 6293 2150
rect 8918 2202 8974 2204
rect 8998 2202 9054 2204
rect 9078 2202 9134 2204
rect 9158 2202 9214 2204
rect 8918 2150 8964 2202
rect 8964 2150 8974 2202
rect 8998 2150 9028 2202
rect 9028 2150 9040 2202
rect 9040 2150 9054 2202
rect 9078 2150 9092 2202
rect 9092 2150 9104 2202
rect 9104 2150 9134 2202
rect 9158 2150 9168 2202
rect 9168 2150 9214 2202
rect 8918 2148 8974 2150
rect 8998 2148 9054 2150
rect 9078 2148 9134 2150
rect 9158 2148 9214 2150
rect 11839 2202 11895 2204
rect 11919 2202 11975 2204
rect 11999 2202 12055 2204
rect 12079 2202 12135 2204
rect 11839 2150 11885 2202
rect 11885 2150 11895 2202
rect 11919 2150 11949 2202
rect 11949 2150 11961 2202
rect 11961 2150 11975 2202
rect 11999 2150 12013 2202
rect 12013 2150 12025 2202
rect 12025 2150 12055 2202
rect 12079 2150 12089 2202
rect 12089 2150 12135 2202
rect 11839 2148 11895 2150
rect 11919 2148 11975 2150
rect 11999 2148 12055 2150
rect 12079 2148 12135 2150
rect 12806 720 12862 776
<< metal3 >>
rect 0 15058 800 15088
rect 4061 15058 4127 15061
rect 0 15056 4127 15058
rect 0 15000 4066 15056
rect 4122 15000 4127 15056
rect 0 14998 4127 15000
rect 0 14968 800 14998
rect 4061 14995 4127 14998
rect 2406 13632 2722 13633
rect 2406 13568 2412 13632
rect 2476 13568 2492 13632
rect 2556 13568 2572 13632
rect 2636 13568 2652 13632
rect 2716 13568 2722 13632
rect 2406 13567 2722 13568
rect 5327 13632 5643 13633
rect 5327 13568 5333 13632
rect 5397 13568 5413 13632
rect 5477 13568 5493 13632
rect 5557 13568 5573 13632
rect 5637 13568 5643 13632
rect 5327 13567 5643 13568
rect 8248 13632 8564 13633
rect 8248 13568 8254 13632
rect 8318 13568 8334 13632
rect 8398 13568 8414 13632
rect 8478 13568 8494 13632
rect 8558 13568 8564 13632
rect 8248 13567 8564 13568
rect 11169 13632 11485 13633
rect 11169 13568 11175 13632
rect 11239 13568 11255 13632
rect 11319 13568 11335 13632
rect 11399 13568 11415 13632
rect 11479 13568 11485 13632
rect 11169 13567 11485 13568
rect 3066 13088 3382 13089
rect 3066 13024 3072 13088
rect 3136 13024 3152 13088
rect 3216 13024 3232 13088
rect 3296 13024 3312 13088
rect 3376 13024 3382 13088
rect 3066 13023 3382 13024
rect 5987 13088 6303 13089
rect 5987 13024 5993 13088
rect 6057 13024 6073 13088
rect 6137 13024 6153 13088
rect 6217 13024 6233 13088
rect 6297 13024 6303 13088
rect 5987 13023 6303 13024
rect 8908 13088 9224 13089
rect 8908 13024 8914 13088
rect 8978 13024 8994 13088
rect 9058 13024 9074 13088
rect 9138 13024 9154 13088
rect 9218 13024 9224 13088
rect 8908 13023 9224 13024
rect 11829 13088 12145 13089
rect 11829 13024 11835 13088
rect 11899 13024 11915 13088
rect 11979 13024 11995 13088
rect 12059 13024 12075 13088
rect 12139 13024 12145 13088
rect 11829 13023 12145 13024
rect 2406 12544 2722 12545
rect 2406 12480 2412 12544
rect 2476 12480 2492 12544
rect 2556 12480 2572 12544
rect 2636 12480 2652 12544
rect 2716 12480 2722 12544
rect 2406 12479 2722 12480
rect 5327 12544 5643 12545
rect 5327 12480 5333 12544
rect 5397 12480 5413 12544
rect 5477 12480 5493 12544
rect 5557 12480 5573 12544
rect 5637 12480 5643 12544
rect 5327 12479 5643 12480
rect 8248 12544 8564 12545
rect 8248 12480 8254 12544
rect 8318 12480 8334 12544
rect 8398 12480 8414 12544
rect 8478 12480 8494 12544
rect 8558 12480 8564 12544
rect 8248 12479 8564 12480
rect 11169 12544 11485 12545
rect 11169 12480 11175 12544
rect 11239 12480 11255 12544
rect 11319 12480 11335 12544
rect 11399 12480 11415 12544
rect 11479 12480 11485 12544
rect 11169 12479 11485 12480
rect 3066 12000 3382 12001
rect 3066 11936 3072 12000
rect 3136 11936 3152 12000
rect 3216 11936 3232 12000
rect 3296 11936 3312 12000
rect 3376 11936 3382 12000
rect 3066 11935 3382 11936
rect 5987 12000 6303 12001
rect 5987 11936 5993 12000
rect 6057 11936 6073 12000
rect 6137 11936 6153 12000
rect 6217 11936 6233 12000
rect 6297 11936 6303 12000
rect 5987 11935 6303 11936
rect 8908 12000 9224 12001
rect 8908 11936 8914 12000
rect 8978 11936 8994 12000
rect 9058 11936 9074 12000
rect 9138 11936 9154 12000
rect 9218 11936 9224 12000
rect 8908 11935 9224 11936
rect 11829 12000 12145 12001
rect 11829 11936 11835 12000
rect 11899 11936 11915 12000
rect 11979 11936 11995 12000
rect 12059 11936 12075 12000
rect 12139 11936 12145 12000
rect 11829 11935 12145 11936
rect 2406 11456 2722 11457
rect 2406 11392 2412 11456
rect 2476 11392 2492 11456
rect 2556 11392 2572 11456
rect 2636 11392 2652 11456
rect 2716 11392 2722 11456
rect 2406 11391 2722 11392
rect 5327 11456 5643 11457
rect 5327 11392 5333 11456
rect 5397 11392 5413 11456
rect 5477 11392 5493 11456
rect 5557 11392 5573 11456
rect 5637 11392 5643 11456
rect 5327 11391 5643 11392
rect 8248 11456 8564 11457
rect 8248 11392 8254 11456
rect 8318 11392 8334 11456
rect 8398 11392 8414 11456
rect 8478 11392 8494 11456
rect 8558 11392 8564 11456
rect 8248 11391 8564 11392
rect 11169 11456 11485 11457
rect 11169 11392 11175 11456
rect 11239 11392 11255 11456
rect 11319 11392 11335 11456
rect 11399 11392 11415 11456
rect 11479 11392 11485 11456
rect 11169 11391 11485 11392
rect 3066 10912 3382 10913
rect 3066 10848 3072 10912
rect 3136 10848 3152 10912
rect 3216 10848 3232 10912
rect 3296 10848 3312 10912
rect 3376 10848 3382 10912
rect 3066 10847 3382 10848
rect 5987 10912 6303 10913
rect 5987 10848 5993 10912
rect 6057 10848 6073 10912
rect 6137 10848 6153 10912
rect 6217 10848 6233 10912
rect 6297 10848 6303 10912
rect 5987 10847 6303 10848
rect 8908 10912 9224 10913
rect 8908 10848 8914 10912
rect 8978 10848 8994 10912
rect 9058 10848 9074 10912
rect 9138 10848 9154 10912
rect 9218 10848 9224 10912
rect 8908 10847 9224 10848
rect 11829 10912 12145 10913
rect 11829 10848 11835 10912
rect 11899 10848 11915 10912
rect 11979 10848 11995 10912
rect 12059 10848 12075 10912
rect 12139 10848 12145 10912
rect 11829 10847 12145 10848
rect 2406 10368 2722 10369
rect 2406 10304 2412 10368
rect 2476 10304 2492 10368
rect 2556 10304 2572 10368
rect 2636 10304 2652 10368
rect 2716 10304 2722 10368
rect 2406 10303 2722 10304
rect 5327 10368 5643 10369
rect 5327 10304 5333 10368
rect 5397 10304 5413 10368
rect 5477 10304 5493 10368
rect 5557 10304 5573 10368
rect 5637 10304 5643 10368
rect 5327 10303 5643 10304
rect 8248 10368 8564 10369
rect 8248 10304 8254 10368
rect 8318 10304 8334 10368
rect 8398 10304 8414 10368
rect 8478 10304 8494 10368
rect 8558 10304 8564 10368
rect 8248 10303 8564 10304
rect 11169 10368 11485 10369
rect 11169 10304 11175 10368
rect 11239 10304 11255 10368
rect 11319 10304 11335 10368
rect 11399 10304 11415 10368
rect 11479 10304 11485 10368
rect 11169 10303 11485 10304
rect 3066 9824 3382 9825
rect 3066 9760 3072 9824
rect 3136 9760 3152 9824
rect 3216 9760 3232 9824
rect 3296 9760 3312 9824
rect 3376 9760 3382 9824
rect 3066 9759 3382 9760
rect 5987 9824 6303 9825
rect 5987 9760 5993 9824
rect 6057 9760 6073 9824
rect 6137 9760 6153 9824
rect 6217 9760 6233 9824
rect 6297 9760 6303 9824
rect 5987 9759 6303 9760
rect 8908 9824 9224 9825
rect 8908 9760 8914 9824
rect 8978 9760 8994 9824
rect 9058 9760 9074 9824
rect 9138 9760 9154 9824
rect 9218 9760 9224 9824
rect 8908 9759 9224 9760
rect 11829 9824 12145 9825
rect 11829 9760 11835 9824
rect 11899 9760 11915 9824
rect 11979 9760 11995 9824
rect 12059 9760 12075 9824
rect 12139 9760 12145 9824
rect 11829 9759 12145 9760
rect 2406 9280 2722 9281
rect 2406 9216 2412 9280
rect 2476 9216 2492 9280
rect 2556 9216 2572 9280
rect 2636 9216 2652 9280
rect 2716 9216 2722 9280
rect 2406 9215 2722 9216
rect 5327 9280 5643 9281
rect 5327 9216 5333 9280
rect 5397 9216 5413 9280
rect 5477 9216 5493 9280
rect 5557 9216 5573 9280
rect 5637 9216 5643 9280
rect 5327 9215 5643 9216
rect 8248 9280 8564 9281
rect 8248 9216 8254 9280
rect 8318 9216 8334 9280
rect 8398 9216 8414 9280
rect 8478 9216 8494 9280
rect 8558 9216 8564 9280
rect 8248 9215 8564 9216
rect 11169 9280 11485 9281
rect 11169 9216 11175 9280
rect 11239 9216 11255 9280
rect 11319 9216 11335 9280
rect 11399 9216 11415 9280
rect 11479 9216 11485 9280
rect 11169 9215 11485 9216
rect 3066 8736 3382 8737
rect 3066 8672 3072 8736
rect 3136 8672 3152 8736
rect 3216 8672 3232 8736
rect 3296 8672 3312 8736
rect 3376 8672 3382 8736
rect 3066 8671 3382 8672
rect 5987 8736 6303 8737
rect 5987 8672 5993 8736
rect 6057 8672 6073 8736
rect 6137 8672 6153 8736
rect 6217 8672 6233 8736
rect 6297 8672 6303 8736
rect 5987 8671 6303 8672
rect 8908 8736 9224 8737
rect 8908 8672 8914 8736
rect 8978 8672 8994 8736
rect 9058 8672 9074 8736
rect 9138 8672 9154 8736
rect 9218 8672 9224 8736
rect 8908 8671 9224 8672
rect 11829 8736 12145 8737
rect 11829 8672 11835 8736
rect 11899 8672 11915 8736
rect 11979 8672 11995 8736
rect 12059 8672 12075 8736
rect 12139 8672 12145 8736
rect 11829 8671 12145 8672
rect 2406 8192 2722 8193
rect 2406 8128 2412 8192
rect 2476 8128 2492 8192
rect 2556 8128 2572 8192
rect 2636 8128 2652 8192
rect 2716 8128 2722 8192
rect 2406 8127 2722 8128
rect 5327 8192 5643 8193
rect 5327 8128 5333 8192
rect 5397 8128 5413 8192
rect 5477 8128 5493 8192
rect 5557 8128 5573 8192
rect 5637 8128 5643 8192
rect 5327 8127 5643 8128
rect 8248 8192 8564 8193
rect 8248 8128 8254 8192
rect 8318 8128 8334 8192
rect 8398 8128 8414 8192
rect 8478 8128 8494 8192
rect 8558 8128 8564 8192
rect 8248 8127 8564 8128
rect 11169 8192 11485 8193
rect 11169 8128 11175 8192
rect 11239 8128 11255 8192
rect 11319 8128 11335 8192
rect 11399 8128 11415 8192
rect 11479 8128 11485 8192
rect 11169 8127 11485 8128
rect 3066 7648 3382 7649
rect 3066 7584 3072 7648
rect 3136 7584 3152 7648
rect 3216 7584 3232 7648
rect 3296 7584 3312 7648
rect 3376 7584 3382 7648
rect 3066 7583 3382 7584
rect 5987 7648 6303 7649
rect 5987 7584 5993 7648
rect 6057 7584 6073 7648
rect 6137 7584 6153 7648
rect 6217 7584 6233 7648
rect 6297 7584 6303 7648
rect 5987 7583 6303 7584
rect 8908 7648 9224 7649
rect 8908 7584 8914 7648
rect 8978 7584 8994 7648
rect 9058 7584 9074 7648
rect 9138 7584 9154 7648
rect 9218 7584 9224 7648
rect 8908 7583 9224 7584
rect 11829 7648 12145 7649
rect 11829 7584 11835 7648
rect 11899 7584 11915 7648
rect 11979 7584 11995 7648
rect 12059 7584 12075 7648
rect 12139 7584 12145 7648
rect 11829 7583 12145 7584
rect 2406 7104 2722 7105
rect 2406 7040 2412 7104
rect 2476 7040 2492 7104
rect 2556 7040 2572 7104
rect 2636 7040 2652 7104
rect 2716 7040 2722 7104
rect 2406 7039 2722 7040
rect 5327 7104 5643 7105
rect 5327 7040 5333 7104
rect 5397 7040 5413 7104
rect 5477 7040 5493 7104
rect 5557 7040 5573 7104
rect 5637 7040 5643 7104
rect 5327 7039 5643 7040
rect 8248 7104 8564 7105
rect 8248 7040 8254 7104
rect 8318 7040 8334 7104
rect 8398 7040 8414 7104
rect 8478 7040 8494 7104
rect 8558 7040 8564 7104
rect 8248 7039 8564 7040
rect 11169 7104 11485 7105
rect 11169 7040 11175 7104
rect 11239 7040 11255 7104
rect 11319 7040 11335 7104
rect 11399 7040 11415 7104
rect 11479 7040 11485 7104
rect 11169 7039 11485 7040
rect 3066 6560 3382 6561
rect 3066 6496 3072 6560
rect 3136 6496 3152 6560
rect 3216 6496 3232 6560
rect 3296 6496 3312 6560
rect 3376 6496 3382 6560
rect 3066 6495 3382 6496
rect 5987 6560 6303 6561
rect 5987 6496 5993 6560
rect 6057 6496 6073 6560
rect 6137 6496 6153 6560
rect 6217 6496 6233 6560
rect 6297 6496 6303 6560
rect 5987 6495 6303 6496
rect 8908 6560 9224 6561
rect 8908 6496 8914 6560
rect 8978 6496 8994 6560
rect 9058 6496 9074 6560
rect 9138 6496 9154 6560
rect 9218 6496 9224 6560
rect 8908 6495 9224 6496
rect 11829 6560 12145 6561
rect 11829 6496 11835 6560
rect 11899 6496 11915 6560
rect 11979 6496 11995 6560
rect 12059 6496 12075 6560
rect 12139 6496 12145 6560
rect 11829 6495 12145 6496
rect 8569 6354 8635 6357
rect 9029 6354 9095 6357
rect 8569 6352 9095 6354
rect 8569 6296 8574 6352
rect 8630 6296 9034 6352
rect 9090 6296 9095 6352
rect 8569 6294 9095 6296
rect 8569 6291 8635 6294
rect 9029 6291 9095 6294
rect 3693 6218 3759 6221
rect 6177 6218 6243 6221
rect 3693 6216 6243 6218
rect 3693 6160 3698 6216
rect 3754 6160 6182 6216
rect 6238 6160 6243 6216
rect 3693 6158 6243 6160
rect 3693 6155 3759 6158
rect 6177 6155 6243 6158
rect 7557 6218 7623 6221
rect 8937 6218 9003 6221
rect 7557 6216 9003 6218
rect 7557 6160 7562 6216
rect 7618 6160 8942 6216
rect 8998 6160 9003 6216
rect 7557 6158 9003 6160
rect 7557 6155 7623 6158
rect 8937 6155 9003 6158
rect 9673 6218 9739 6221
rect 10225 6218 10291 6221
rect 9673 6216 10291 6218
rect 9673 6160 9678 6216
rect 9734 6160 10230 6216
rect 10286 6160 10291 6216
rect 9673 6158 10291 6160
rect 9673 6155 9739 6158
rect 10225 6155 10291 6158
rect 2406 6016 2722 6017
rect 2406 5952 2412 6016
rect 2476 5952 2492 6016
rect 2556 5952 2572 6016
rect 2636 5952 2652 6016
rect 2716 5952 2722 6016
rect 2406 5951 2722 5952
rect 5327 6016 5643 6017
rect 5327 5952 5333 6016
rect 5397 5952 5413 6016
rect 5477 5952 5493 6016
rect 5557 5952 5573 6016
rect 5637 5952 5643 6016
rect 5327 5951 5643 5952
rect 8248 6016 8564 6017
rect 8248 5952 8254 6016
rect 8318 5952 8334 6016
rect 8398 5952 8414 6016
rect 8478 5952 8494 6016
rect 8558 5952 8564 6016
rect 8248 5951 8564 5952
rect 11169 6016 11485 6017
rect 11169 5952 11175 6016
rect 11239 5952 11255 6016
rect 11319 5952 11335 6016
rect 11399 5952 11415 6016
rect 11479 5952 11485 6016
rect 11169 5951 11485 5952
rect 7741 5674 7807 5677
rect 9305 5674 9371 5677
rect 7741 5672 9371 5674
rect 7741 5616 7746 5672
rect 7802 5616 9310 5672
rect 9366 5616 9371 5672
rect 7741 5614 9371 5616
rect 7741 5611 7807 5614
rect 9305 5611 9371 5614
rect 3066 5472 3382 5473
rect 3066 5408 3072 5472
rect 3136 5408 3152 5472
rect 3216 5408 3232 5472
rect 3296 5408 3312 5472
rect 3376 5408 3382 5472
rect 3066 5407 3382 5408
rect 5987 5472 6303 5473
rect 5987 5408 5993 5472
rect 6057 5408 6073 5472
rect 6137 5408 6153 5472
rect 6217 5408 6233 5472
rect 6297 5408 6303 5472
rect 5987 5407 6303 5408
rect 8908 5472 9224 5473
rect 8908 5408 8914 5472
rect 8978 5408 8994 5472
rect 9058 5408 9074 5472
rect 9138 5408 9154 5472
rect 9218 5408 9224 5472
rect 8908 5407 9224 5408
rect 11829 5472 12145 5473
rect 11829 5408 11835 5472
rect 11899 5408 11915 5472
rect 11979 5408 11995 5472
rect 12059 5408 12075 5472
rect 12139 5408 12145 5472
rect 11829 5407 12145 5408
rect 4153 5266 4219 5269
rect 6269 5266 6335 5269
rect 6913 5266 6979 5269
rect 4153 5264 6979 5266
rect 4153 5208 4158 5264
rect 4214 5208 6274 5264
rect 6330 5208 6918 5264
rect 6974 5208 6979 5264
rect 4153 5206 6979 5208
rect 4153 5203 4219 5206
rect 6269 5203 6335 5206
rect 6913 5203 6979 5206
rect 3877 5130 3943 5133
rect 7097 5130 7163 5133
rect 8385 5130 8451 5133
rect 3877 5128 8451 5130
rect 3877 5072 3882 5128
rect 3938 5072 7102 5128
rect 7158 5072 8390 5128
rect 8446 5072 8451 5128
rect 3877 5070 8451 5072
rect 3877 5067 3943 5070
rect 7097 5067 7163 5070
rect 8385 5067 8451 5070
rect 2406 4928 2722 4929
rect 2406 4864 2412 4928
rect 2476 4864 2492 4928
rect 2556 4864 2572 4928
rect 2636 4864 2652 4928
rect 2716 4864 2722 4928
rect 2406 4863 2722 4864
rect 5327 4928 5643 4929
rect 5327 4864 5333 4928
rect 5397 4864 5413 4928
rect 5477 4864 5493 4928
rect 5557 4864 5573 4928
rect 5637 4864 5643 4928
rect 5327 4863 5643 4864
rect 8248 4928 8564 4929
rect 8248 4864 8254 4928
rect 8318 4864 8334 4928
rect 8398 4864 8414 4928
rect 8478 4864 8494 4928
rect 8558 4864 8564 4928
rect 8248 4863 8564 4864
rect 11169 4928 11485 4929
rect 11169 4864 11175 4928
rect 11239 4864 11255 4928
rect 11319 4864 11335 4928
rect 11399 4864 11415 4928
rect 11479 4864 11485 4928
rect 11169 4863 11485 4864
rect 8937 4586 9003 4589
rect 8937 4584 9506 4586
rect 8937 4528 8942 4584
rect 8998 4528 9506 4584
rect 8937 4526 9506 4528
rect 8937 4523 9003 4526
rect 3066 4384 3382 4385
rect 3066 4320 3072 4384
rect 3136 4320 3152 4384
rect 3216 4320 3232 4384
rect 3296 4320 3312 4384
rect 3376 4320 3382 4384
rect 3066 4319 3382 4320
rect 5987 4384 6303 4385
rect 5987 4320 5993 4384
rect 6057 4320 6073 4384
rect 6137 4320 6153 4384
rect 6217 4320 6233 4384
rect 6297 4320 6303 4384
rect 5987 4319 6303 4320
rect 8908 4384 9224 4385
rect 8908 4320 8914 4384
rect 8978 4320 8994 4384
rect 9058 4320 9074 4384
rect 9138 4320 9154 4384
rect 9218 4320 9224 4384
rect 8908 4319 9224 4320
rect 9446 4317 9506 4526
rect 11829 4384 12145 4385
rect 11829 4320 11835 4384
rect 11899 4320 11915 4384
rect 11979 4320 11995 4384
rect 12059 4320 12075 4384
rect 12139 4320 12145 4384
rect 11829 4319 12145 4320
rect 9397 4312 9506 4317
rect 9397 4256 9402 4312
rect 9458 4256 9506 4312
rect 9397 4254 9506 4256
rect 9397 4251 9463 4254
rect 1485 4178 1551 4181
rect 3049 4178 3115 4181
rect 1485 4176 3115 4178
rect 1485 4120 1490 4176
rect 1546 4120 3054 4176
rect 3110 4120 3115 4176
rect 1485 4118 3115 4120
rect 1485 4115 1551 4118
rect 3049 4115 3115 4118
rect 5073 4178 5139 4181
rect 5717 4178 5783 4181
rect 7925 4178 7991 4181
rect 5073 4176 7991 4178
rect 5073 4120 5078 4176
rect 5134 4120 5722 4176
rect 5778 4120 7930 4176
rect 7986 4120 7991 4176
rect 5073 4118 7991 4120
rect 5073 4115 5139 4118
rect 5717 4115 5783 4118
rect 7925 4115 7991 4118
rect 2406 3840 2722 3841
rect 2406 3776 2412 3840
rect 2476 3776 2492 3840
rect 2556 3776 2572 3840
rect 2636 3776 2652 3840
rect 2716 3776 2722 3840
rect 2406 3775 2722 3776
rect 5327 3840 5643 3841
rect 5327 3776 5333 3840
rect 5397 3776 5413 3840
rect 5477 3776 5493 3840
rect 5557 3776 5573 3840
rect 5637 3776 5643 3840
rect 5327 3775 5643 3776
rect 8248 3840 8564 3841
rect 8248 3776 8254 3840
rect 8318 3776 8334 3840
rect 8398 3776 8414 3840
rect 8478 3776 8494 3840
rect 8558 3776 8564 3840
rect 8248 3775 8564 3776
rect 11169 3840 11485 3841
rect 11169 3776 11175 3840
rect 11239 3776 11255 3840
rect 11319 3776 11335 3840
rect 11399 3776 11415 3840
rect 11479 3776 11485 3840
rect 11169 3775 11485 3776
rect 4981 3634 5047 3637
rect 7005 3634 7071 3637
rect 4981 3632 7071 3634
rect 4981 3576 4986 3632
rect 5042 3576 7010 3632
rect 7066 3576 7071 3632
rect 4981 3574 7071 3576
rect 4981 3571 5047 3574
rect 7005 3571 7071 3574
rect 4705 3498 4771 3501
rect 7925 3498 7991 3501
rect 4705 3496 7991 3498
rect 4705 3440 4710 3496
rect 4766 3440 7930 3496
rect 7986 3440 7991 3496
rect 4705 3438 7991 3440
rect 4705 3435 4771 3438
rect 7925 3435 7991 3438
rect 3066 3296 3382 3297
rect 3066 3232 3072 3296
rect 3136 3232 3152 3296
rect 3216 3232 3232 3296
rect 3296 3232 3312 3296
rect 3376 3232 3382 3296
rect 3066 3231 3382 3232
rect 5987 3296 6303 3297
rect 5987 3232 5993 3296
rect 6057 3232 6073 3296
rect 6137 3232 6153 3296
rect 6217 3232 6233 3296
rect 6297 3232 6303 3296
rect 5987 3231 6303 3232
rect 8908 3296 9224 3297
rect 8908 3232 8914 3296
rect 8978 3232 8994 3296
rect 9058 3232 9074 3296
rect 9138 3232 9154 3296
rect 9218 3232 9224 3296
rect 8908 3231 9224 3232
rect 11829 3296 12145 3297
rect 11829 3232 11835 3296
rect 11899 3232 11915 3296
rect 11979 3232 11995 3296
rect 12059 3232 12075 3296
rect 12139 3232 12145 3296
rect 11829 3231 12145 3232
rect 1577 3090 1643 3093
rect 4429 3090 4495 3093
rect 1577 3088 4495 3090
rect 1577 3032 1582 3088
rect 1638 3032 4434 3088
rect 4490 3032 4495 3088
rect 1577 3030 4495 3032
rect 1577 3027 1643 3030
rect 4429 3027 4495 3030
rect 4889 2954 4955 2957
rect 9029 2954 9095 2957
rect 4889 2952 9095 2954
rect 4889 2896 4894 2952
rect 4950 2896 9034 2952
rect 9090 2896 9095 2952
rect 4889 2894 9095 2896
rect 4889 2891 4955 2894
rect 9029 2891 9095 2894
rect 4153 2818 4219 2821
rect 5073 2818 5139 2821
rect 4153 2816 5139 2818
rect 4153 2760 4158 2816
rect 4214 2760 5078 2816
rect 5134 2760 5139 2816
rect 4153 2758 5139 2760
rect 4153 2755 4219 2758
rect 5073 2755 5139 2758
rect 2406 2752 2722 2753
rect 2406 2688 2412 2752
rect 2476 2688 2492 2752
rect 2556 2688 2572 2752
rect 2636 2688 2652 2752
rect 2716 2688 2722 2752
rect 2406 2687 2722 2688
rect 5327 2752 5643 2753
rect 5327 2688 5333 2752
rect 5397 2688 5413 2752
rect 5477 2688 5493 2752
rect 5557 2688 5573 2752
rect 5637 2688 5643 2752
rect 5327 2687 5643 2688
rect 8248 2752 8564 2753
rect 8248 2688 8254 2752
rect 8318 2688 8334 2752
rect 8398 2688 8414 2752
rect 8478 2688 8494 2752
rect 8558 2688 8564 2752
rect 8248 2687 8564 2688
rect 11169 2752 11485 2753
rect 11169 2688 11175 2752
rect 11239 2688 11255 2752
rect 11319 2688 11335 2752
rect 11399 2688 11415 2752
rect 11479 2688 11485 2752
rect 11169 2687 11485 2688
rect 3066 2208 3382 2209
rect 3066 2144 3072 2208
rect 3136 2144 3152 2208
rect 3216 2144 3232 2208
rect 3296 2144 3312 2208
rect 3376 2144 3382 2208
rect 3066 2143 3382 2144
rect 5987 2208 6303 2209
rect 5987 2144 5993 2208
rect 6057 2144 6073 2208
rect 6137 2144 6153 2208
rect 6217 2144 6233 2208
rect 6297 2144 6303 2208
rect 5987 2143 6303 2144
rect 8908 2208 9224 2209
rect 8908 2144 8914 2208
rect 8978 2144 8994 2208
rect 9058 2144 9074 2208
rect 9138 2144 9154 2208
rect 9218 2144 9224 2208
rect 8908 2143 9224 2144
rect 11829 2208 12145 2209
rect 11829 2144 11835 2208
rect 11899 2144 11915 2208
rect 11979 2144 11995 2208
rect 12059 2144 12075 2208
rect 12139 2144 12145 2208
rect 11829 2143 12145 2144
rect 12801 778 12867 781
rect 13122 778 13922 808
rect 12801 776 13922 778
rect 12801 720 12806 776
rect 12862 720 13922 776
rect 12801 718 13922 720
rect 12801 715 12867 718
rect 13122 688 13922 718
<< via3 >>
rect 2412 13628 2476 13632
rect 2412 13572 2416 13628
rect 2416 13572 2472 13628
rect 2472 13572 2476 13628
rect 2412 13568 2476 13572
rect 2492 13628 2556 13632
rect 2492 13572 2496 13628
rect 2496 13572 2552 13628
rect 2552 13572 2556 13628
rect 2492 13568 2556 13572
rect 2572 13628 2636 13632
rect 2572 13572 2576 13628
rect 2576 13572 2632 13628
rect 2632 13572 2636 13628
rect 2572 13568 2636 13572
rect 2652 13628 2716 13632
rect 2652 13572 2656 13628
rect 2656 13572 2712 13628
rect 2712 13572 2716 13628
rect 2652 13568 2716 13572
rect 5333 13628 5397 13632
rect 5333 13572 5337 13628
rect 5337 13572 5393 13628
rect 5393 13572 5397 13628
rect 5333 13568 5397 13572
rect 5413 13628 5477 13632
rect 5413 13572 5417 13628
rect 5417 13572 5473 13628
rect 5473 13572 5477 13628
rect 5413 13568 5477 13572
rect 5493 13628 5557 13632
rect 5493 13572 5497 13628
rect 5497 13572 5553 13628
rect 5553 13572 5557 13628
rect 5493 13568 5557 13572
rect 5573 13628 5637 13632
rect 5573 13572 5577 13628
rect 5577 13572 5633 13628
rect 5633 13572 5637 13628
rect 5573 13568 5637 13572
rect 8254 13628 8318 13632
rect 8254 13572 8258 13628
rect 8258 13572 8314 13628
rect 8314 13572 8318 13628
rect 8254 13568 8318 13572
rect 8334 13628 8398 13632
rect 8334 13572 8338 13628
rect 8338 13572 8394 13628
rect 8394 13572 8398 13628
rect 8334 13568 8398 13572
rect 8414 13628 8478 13632
rect 8414 13572 8418 13628
rect 8418 13572 8474 13628
rect 8474 13572 8478 13628
rect 8414 13568 8478 13572
rect 8494 13628 8558 13632
rect 8494 13572 8498 13628
rect 8498 13572 8554 13628
rect 8554 13572 8558 13628
rect 8494 13568 8558 13572
rect 11175 13628 11239 13632
rect 11175 13572 11179 13628
rect 11179 13572 11235 13628
rect 11235 13572 11239 13628
rect 11175 13568 11239 13572
rect 11255 13628 11319 13632
rect 11255 13572 11259 13628
rect 11259 13572 11315 13628
rect 11315 13572 11319 13628
rect 11255 13568 11319 13572
rect 11335 13628 11399 13632
rect 11335 13572 11339 13628
rect 11339 13572 11395 13628
rect 11395 13572 11399 13628
rect 11335 13568 11399 13572
rect 11415 13628 11479 13632
rect 11415 13572 11419 13628
rect 11419 13572 11475 13628
rect 11475 13572 11479 13628
rect 11415 13568 11479 13572
rect 3072 13084 3136 13088
rect 3072 13028 3076 13084
rect 3076 13028 3132 13084
rect 3132 13028 3136 13084
rect 3072 13024 3136 13028
rect 3152 13084 3216 13088
rect 3152 13028 3156 13084
rect 3156 13028 3212 13084
rect 3212 13028 3216 13084
rect 3152 13024 3216 13028
rect 3232 13084 3296 13088
rect 3232 13028 3236 13084
rect 3236 13028 3292 13084
rect 3292 13028 3296 13084
rect 3232 13024 3296 13028
rect 3312 13084 3376 13088
rect 3312 13028 3316 13084
rect 3316 13028 3372 13084
rect 3372 13028 3376 13084
rect 3312 13024 3376 13028
rect 5993 13084 6057 13088
rect 5993 13028 5997 13084
rect 5997 13028 6053 13084
rect 6053 13028 6057 13084
rect 5993 13024 6057 13028
rect 6073 13084 6137 13088
rect 6073 13028 6077 13084
rect 6077 13028 6133 13084
rect 6133 13028 6137 13084
rect 6073 13024 6137 13028
rect 6153 13084 6217 13088
rect 6153 13028 6157 13084
rect 6157 13028 6213 13084
rect 6213 13028 6217 13084
rect 6153 13024 6217 13028
rect 6233 13084 6297 13088
rect 6233 13028 6237 13084
rect 6237 13028 6293 13084
rect 6293 13028 6297 13084
rect 6233 13024 6297 13028
rect 8914 13084 8978 13088
rect 8914 13028 8918 13084
rect 8918 13028 8974 13084
rect 8974 13028 8978 13084
rect 8914 13024 8978 13028
rect 8994 13084 9058 13088
rect 8994 13028 8998 13084
rect 8998 13028 9054 13084
rect 9054 13028 9058 13084
rect 8994 13024 9058 13028
rect 9074 13084 9138 13088
rect 9074 13028 9078 13084
rect 9078 13028 9134 13084
rect 9134 13028 9138 13084
rect 9074 13024 9138 13028
rect 9154 13084 9218 13088
rect 9154 13028 9158 13084
rect 9158 13028 9214 13084
rect 9214 13028 9218 13084
rect 9154 13024 9218 13028
rect 11835 13084 11899 13088
rect 11835 13028 11839 13084
rect 11839 13028 11895 13084
rect 11895 13028 11899 13084
rect 11835 13024 11899 13028
rect 11915 13084 11979 13088
rect 11915 13028 11919 13084
rect 11919 13028 11975 13084
rect 11975 13028 11979 13084
rect 11915 13024 11979 13028
rect 11995 13084 12059 13088
rect 11995 13028 11999 13084
rect 11999 13028 12055 13084
rect 12055 13028 12059 13084
rect 11995 13024 12059 13028
rect 12075 13084 12139 13088
rect 12075 13028 12079 13084
rect 12079 13028 12135 13084
rect 12135 13028 12139 13084
rect 12075 13024 12139 13028
rect 2412 12540 2476 12544
rect 2412 12484 2416 12540
rect 2416 12484 2472 12540
rect 2472 12484 2476 12540
rect 2412 12480 2476 12484
rect 2492 12540 2556 12544
rect 2492 12484 2496 12540
rect 2496 12484 2552 12540
rect 2552 12484 2556 12540
rect 2492 12480 2556 12484
rect 2572 12540 2636 12544
rect 2572 12484 2576 12540
rect 2576 12484 2632 12540
rect 2632 12484 2636 12540
rect 2572 12480 2636 12484
rect 2652 12540 2716 12544
rect 2652 12484 2656 12540
rect 2656 12484 2712 12540
rect 2712 12484 2716 12540
rect 2652 12480 2716 12484
rect 5333 12540 5397 12544
rect 5333 12484 5337 12540
rect 5337 12484 5393 12540
rect 5393 12484 5397 12540
rect 5333 12480 5397 12484
rect 5413 12540 5477 12544
rect 5413 12484 5417 12540
rect 5417 12484 5473 12540
rect 5473 12484 5477 12540
rect 5413 12480 5477 12484
rect 5493 12540 5557 12544
rect 5493 12484 5497 12540
rect 5497 12484 5553 12540
rect 5553 12484 5557 12540
rect 5493 12480 5557 12484
rect 5573 12540 5637 12544
rect 5573 12484 5577 12540
rect 5577 12484 5633 12540
rect 5633 12484 5637 12540
rect 5573 12480 5637 12484
rect 8254 12540 8318 12544
rect 8254 12484 8258 12540
rect 8258 12484 8314 12540
rect 8314 12484 8318 12540
rect 8254 12480 8318 12484
rect 8334 12540 8398 12544
rect 8334 12484 8338 12540
rect 8338 12484 8394 12540
rect 8394 12484 8398 12540
rect 8334 12480 8398 12484
rect 8414 12540 8478 12544
rect 8414 12484 8418 12540
rect 8418 12484 8474 12540
rect 8474 12484 8478 12540
rect 8414 12480 8478 12484
rect 8494 12540 8558 12544
rect 8494 12484 8498 12540
rect 8498 12484 8554 12540
rect 8554 12484 8558 12540
rect 8494 12480 8558 12484
rect 11175 12540 11239 12544
rect 11175 12484 11179 12540
rect 11179 12484 11235 12540
rect 11235 12484 11239 12540
rect 11175 12480 11239 12484
rect 11255 12540 11319 12544
rect 11255 12484 11259 12540
rect 11259 12484 11315 12540
rect 11315 12484 11319 12540
rect 11255 12480 11319 12484
rect 11335 12540 11399 12544
rect 11335 12484 11339 12540
rect 11339 12484 11395 12540
rect 11395 12484 11399 12540
rect 11335 12480 11399 12484
rect 11415 12540 11479 12544
rect 11415 12484 11419 12540
rect 11419 12484 11475 12540
rect 11475 12484 11479 12540
rect 11415 12480 11479 12484
rect 3072 11996 3136 12000
rect 3072 11940 3076 11996
rect 3076 11940 3132 11996
rect 3132 11940 3136 11996
rect 3072 11936 3136 11940
rect 3152 11996 3216 12000
rect 3152 11940 3156 11996
rect 3156 11940 3212 11996
rect 3212 11940 3216 11996
rect 3152 11936 3216 11940
rect 3232 11996 3296 12000
rect 3232 11940 3236 11996
rect 3236 11940 3292 11996
rect 3292 11940 3296 11996
rect 3232 11936 3296 11940
rect 3312 11996 3376 12000
rect 3312 11940 3316 11996
rect 3316 11940 3372 11996
rect 3372 11940 3376 11996
rect 3312 11936 3376 11940
rect 5993 11996 6057 12000
rect 5993 11940 5997 11996
rect 5997 11940 6053 11996
rect 6053 11940 6057 11996
rect 5993 11936 6057 11940
rect 6073 11996 6137 12000
rect 6073 11940 6077 11996
rect 6077 11940 6133 11996
rect 6133 11940 6137 11996
rect 6073 11936 6137 11940
rect 6153 11996 6217 12000
rect 6153 11940 6157 11996
rect 6157 11940 6213 11996
rect 6213 11940 6217 11996
rect 6153 11936 6217 11940
rect 6233 11996 6297 12000
rect 6233 11940 6237 11996
rect 6237 11940 6293 11996
rect 6293 11940 6297 11996
rect 6233 11936 6297 11940
rect 8914 11996 8978 12000
rect 8914 11940 8918 11996
rect 8918 11940 8974 11996
rect 8974 11940 8978 11996
rect 8914 11936 8978 11940
rect 8994 11996 9058 12000
rect 8994 11940 8998 11996
rect 8998 11940 9054 11996
rect 9054 11940 9058 11996
rect 8994 11936 9058 11940
rect 9074 11996 9138 12000
rect 9074 11940 9078 11996
rect 9078 11940 9134 11996
rect 9134 11940 9138 11996
rect 9074 11936 9138 11940
rect 9154 11996 9218 12000
rect 9154 11940 9158 11996
rect 9158 11940 9214 11996
rect 9214 11940 9218 11996
rect 9154 11936 9218 11940
rect 11835 11996 11899 12000
rect 11835 11940 11839 11996
rect 11839 11940 11895 11996
rect 11895 11940 11899 11996
rect 11835 11936 11899 11940
rect 11915 11996 11979 12000
rect 11915 11940 11919 11996
rect 11919 11940 11975 11996
rect 11975 11940 11979 11996
rect 11915 11936 11979 11940
rect 11995 11996 12059 12000
rect 11995 11940 11999 11996
rect 11999 11940 12055 11996
rect 12055 11940 12059 11996
rect 11995 11936 12059 11940
rect 12075 11996 12139 12000
rect 12075 11940 12079 11996
rect 12079 11940 12135 11996
rect 12135 11940 12139 11996
rect 12075 11936 12139 11940
rect 2412 11452 2476 11456
rect 2412 11396 2416 11452
rect 2416 11396 2472 11452
rect 2472 11396 2476 11452
rect 2412 11392 2476 11396
rect 2492 11452 2556 11456
rect 2492 11396 2496 11452
rect 2496 11396 2552 11452
rect 2552 11396 2556 11452
rect 2492 11392 2556 11396
rect 2572 11452 2636 11456
rect 2572 11396 2576 11452
rect 2576 11396 2632 11452
rect 2632 11396 2636 11452
rect 2572 11392 2636 11396
rect 2652 11452 2716 11456
rect 2652 11396 2656 11452
rect 2656 11396 2712 11452
rect 2712 11396 2716 11452
rect 2652 11392 2716 11396
rect 5333 11452 5397 11456
rect 5333 11396 5337 11452
rect 5337 11396 5393 11452
rect 5393 11396 5397 11452
rect 5333 11392 5397 11396
rect 5413 11452 5477 11456
rect 5413 11396 5417 11452
rect 5417 11396 5473 11452
rect 5473 11396 5477 11452
rect 5413 11392 5477 11396
rect 5493 11452 5557 11456
rect 5493 11396 5497 11452
rect 5497 11396 5553 11452
rect 5553 11396 5557 11452
rect 5493 11392 5557 11396
rect 5573 11452 5637 11456
rect 5573 11396 5577 11452
rect 5577 11396 5633 11452
rect 5633 11396 5637 11452
rect 5573 11392 5637 11396
rect 8254 11452 8318 11456
rect 8254 11396 8258 11452
rect 8258 11396 8314 11452
rect 8314 11396 8318 11452
rect 8254 11392 8318 11396
rect 8334 11452 8398 11456
rect 8334 11396 8338 11452
rect 8338 11396 8394 11452
rect 8394 11396 8398 11452
rect 8334 11392 8398 11396
rect 8414 11452 8478 11456
rect 8414 11396 8418 11452
rect 8418 11396 8474 11452
rect 8474 11396 8478 11452
rect 8414 11392 8478 11396
rect 8494 11452 8558 11456
rect 8494 11396 8498 11452
rect 8498 11396 8554 11452
rect 8554 11396 8558 11452
rect 8494 11392 8558 11396
rect 11175 11452 11239 11456
rect 11175 11396 11179 11452
rect 11179 11396 11235 11452
rect 11235 11396 11239 11452
rect 11175 11392 11239 11396
rect 11255 11452 11319 11456
rect 11255 11396 11259 11452
rect 11259 11396 11315 11452
rect 11315 11396 11319 11452
rect 11255 11392 11319 11396
rect 11335 11452 11399 11456
rect 11335 11396 11339 11452
rect 11339 11396 11395 11452
rect 11395 11396 11399 11452
rect 11335 11392 11399 11396
rect 11415 11452 11479 11456
rect 11415 11396 11419 11452
rect 11419 11396 11475 11452
rect 11475 11396 11479 11452
rect 11415 11392 11479 11396
rect 3072 10908 3136 10912
rect 3072 10852 3076 10908
rect 3076 10852 3132 10908
rect 3132 10852 3136 10908
rect 3072 10848 3136 10852
rect 3152 10908 3216 10912
rect 3152 10852 3156 10908
rect 3156 10852 3212 10908
rect 3212 10852 3216 10908
rect 3152 10848 3216 10852
rect 3232 10908 3296 10912
rect 3232 10852 3236 10908
rect 3236 10852 3292 10908
rect 3292 10852 3296 10908
rect 3232 10848 3296 10852
rect 3312 10908 3376 10912
rect 3312 10852 3316 10908
rect 3316 10852 3372 10908
rect 3372 10852 3376 10908
rect 3312 10848 3376 10852
rect 5993 10908 6057 10912
rect 5993 10852 5997 10908
rect 5997 10852 6053 10908
rect 6053 10852 6057 10908
rect 5993 10848 6057 10852
rect 6073 10908 6137 10912
rect 6073 10852 6077 10908
rect 6077 10852 6133 10908
rect 6133 10852 6137 10908
rect 6073 10848 6137 10852
rect 6153 10908 6217 10912
rect 6153 10852 6157 10908
rect 6157 10852 6213 10908
rect 6213 10852 6217 10908
rect 6153 10848 6217 10852
rect 6233 10908 6297 10912
rect 6233 10852 6237 10908
rect 6237 10852 6293 10908
rect 6293 10852 6297 10908
rect 6233 10848 6297 10852
rect 8914 10908 8978 10912
rect 8914 10852 8918 10908
rect 8918 10852 8974 10908
rect 8974 10852 8978 10908
rect 8914 10848 8978 10852
rect 8994 10908 9058 10912
rect 8994 10852 8998 10908
rect 8998 10852 9054 10908
rect 9054 10852 9058 10908
rect 8994 10848 9058 10852
rect 9074 10908 9138 10912
rect 9074 10852 9078 10908
rect 9078 10852 9134 10908
rect 9134 10852 9138 10908
rect 9074 10848 9138 10852
rect 9154 10908 9218 10912
rect 9154 10852 9158 10908
rect 9158 10852 9214 10908
rect 9214 10852 9218 10908
rect 9154 10848 9218 10852
rect 11835 10908 11899 10912
rect 11835 10852 11839 10908
rect 11839 10852 11895 10908
rect 11895 10852 11899 10908
rect 11835 10848 11899 10852
rect 11915 10908 11979 10912
rect 11915 10852 11919 10908
rect 11919 10852 11975 10908
rect 11975 10852 11979 10908
rect 11915 10848 11979 10852
rect 11995 10908 12059 10912
rect 11995 10852 11999 10908
rect 11999 10852 12055 10908
rect 12055 10852 12059 10908
rect 11995 10848 12059 10852
rect 12075 10908 12139 10912
rect 12075 10852 12079 10908
rect 12079 10852 12135 10908
rect 12135 10852 12139 10908
rect 12075 10848 12139 10852
rect 2412 10364 2476 10368
rect 2412 10308 2416 10364
rect 2416 10308 2472 10364
rect 2472 10308 2476 10364
rect 2412 10304 2476 10308
rect 2492 10364 2556 10368
rect 2492 10308 2496 10364
rect 2496 10308 2552 10364
rect 2552 10308 2556 10364
rect 2492 10304 2556 10308
rect 2572 10364 2636 10368
rect 2572 10308 2576 10364
rect 2576 10308 2632 10364
rect 2632 10308 2636 10364
rect 2572 10304 2636 10308
rect 2652 10364 2716 10368
rect 2652 10308 2656 10364
rect 2656 10308 2712 10364
rect 2712 10308 2716 10364
rect 2652 10304 2716 10308
rect 5333 10364 5397 10368
rect 5333 10308 5337 10364
rect 5337 10308 5393 10364
rect 5393 10308 5397 10364
rect 5333 10304 5397 10308
rect 5413 10364 5477 10368
rect 5413 10308 5417 10364
rect 5417 10308 5473 10364
rect 5473 10308 5477 10364
rect 5413 10304 5477 10308
rect 5493 10364 5557 10368
rect 5493 10308 5497 10364
rect 5497 10308 5553 10364
rect 5553 10308 5557 10364
rect 5493 10304 5557 10308
rect 5573 10364 5637 10368
rect 5573 10308 5577 10364
rect 5577 10308 5633 10364
rect 5633 10308 5637 10364
rect 5573 10304 5637 10308
rect 8254 10364 8318 10368
rect 8254 10308 8258 10364
rect 8258 10308 8314 10364
rect 8314 10308 8318 10364
rect 8254 10304 8318 10308
rect 8334 10364 8398 10368
rect 8334 10308 8338 10364
rect 8338 10308 8394 10364
rect 8394 10308 8398 10364
rect 8334 10304 8398 10308
rect 8414 10364 8478 10368
rect 8414 10308 8418 10364
rect 8418 10308 8474 10364
rect 8474 10308 8478 10364
rect 8414 10304 8478 10308
rect 8494 10364 8558 10368
rect 8494 10308 8498 10364
rect 8498 10308 8554 10364
rect 8554 10308 8558 10364
rect 8494 10304 8558 10308
rect 11175 10364 11239 10368
rect 11175 10308 11179 10364
rect 11179 10308 11235 10364
rect 11235 10308 11239 10364
rect 11175 10304 11239 10308
rect 11255 10364 11319 10368
rect 11255 10308 11259 10364
rect 11259 10308 11315 10364
rect 11315 10308 11319 10364
rect 11255 10304 11319 10308
rect 11335 10364 11399 10368
rect 11335 10308 11339 10364
rect 11339 10308 11395 10364
rect 11395 10308 11399 10364
rect 11335 10304 11399 10308
rect 11415 10364 11479 10368
rect 11415 10308 11419 10364
rect 11419 10308 11475 10364
rect 11475 10308 11479 10364
rect 11415 10304 11479 10308
rect 3072 9820 3136 9824
rect 3072 9764 3076 9820
rect 3076 9764 3132 9820
rect 3132 9764 3136 9820
rect 3072 9760 3136 9764
rect 3152 9820 3216 9824
rect 3152 9764 3156 9820
rect 3156 9764 3212 9820
rect 3212 9764 3216 9820
rect 3152 9760 3216 9764
rect 3232 9820 3296 9824
rect 3232 9764 3236 9820
rect 3236 9764 3292 9820
rect 3292 9764 3296 9820
rect 3232 9760 3296 9764
rect 3312 9820 3376 9824
rect 3312 9764 3316 9820
rect 3316 9764 3372 9820
rect 3372 9764 3376 9820
rect 3312 9760 3376 9764
rect 5993 9820 6057 9824
rect 5993 9764 5997 9820
rect 5997 9764 6053 9820
rect 6053 9764 6057 9820
rect 5993 9760 6057 9764
rect 6073 9820 6137 9824
rect 6073 9764 6077 9820
rect 6077 9764 6133 9820
rect 6133 9764 6137 9820
rect 6073 9760 6137 9764
rect 6153 9820 6217 9824
rect 6153 9764 6157 9820
rect 6157 9764 6213 9820
rect 6213 9764 6217 9820
rect 6153 9760 6217 9764
rect 6233 9820 6297 9824
rect 6233 9764 6237 9820
rect 6237 9764 6293 9820
rect 6293 9764 6297 9820
rect 6233 9760 6297 9764
rect 8914 9820 8978 9824
rect 8914 9764 8918 9820
rect 8918 9764 8974 9820
rect 8974 9764 8978 9820
rect 8914 9760 8978 9764
rect 8994 9820 9058 9824
rect 8994 9764 8998 9820
rect 8998 9764 9054 9820
rect 9054 9764 9058 9820
rect 8994 9760 9058 9764
rect 9074 9820 9138 9824
rect 9074 9764 9078 9820
rect 9078 9764 9134 9820
rect 9134 9764 9138 9820
rect 9074 9760 9138 9764
rect 9154 9820 9218 9824
rect 9154 9764 9158 9820
rect 9158 9764 9214 9820
rect 9214 9764 9218 9820
rect 9154 9760 9218 9764
rect 11835 9820 11899 9824
rect 11835 9764 11839 9820
rect 11839 9764 11895 9820
rect 11895 9764 11899 9820
rect 11835 9760 11899 9764
rect 11915 9820 11979 9824
rect 11915 9764 11919 9820
rect 11919 9764 11975 9820
rect 11975 9764 11979 9820
rect 11915 9760 11979 9764
rect 11995 9820 12059 9824
rect 11995 9764 11999 9820
rect 11999 9764 12055 9820
rect 12055 9764 12059 9820
rect 11995 9760 12059 9764
rect 12075 9820 12139 9824
rect 12075 9764 12079 9820
rect 12079 9764 12135 9820
rect 12135 9764 12139 9820
rect 12075 9760 12139 9764
rect 2412 9276 2476 9280
rect 2412 9220 2416 9276
rect 2416 9220 2472 9276
rect 2472 9220 2476 9276
rect 2412 9216 2476 9220
rect 2492 9276 2556 9280
rect 2492 9220 2496 9276
rect 2496 9220 2552 9276
rect 2552 9220 2556 9276
rect 2492 9216 2556 9220
rect 2572 9276 2636 9280
rect 2572 9220 2576 9276
rect 2576 9220 2632 9276
rect 2632 9220 2636 9276
rect 2572 9216 2636 9220
rect 2652 9276 2716 9280
rect 2652 9220 2656 9276
rect 2656 9220 2712 9276
rect 2712 9220 2716 9276
rect 2652 9216 2716 9220
rect 5333 9276 5397 9280
rect 5333 9220 5337 9276
rect 5337 9220 5393 9276
rect 5393 9220 5397 9276
rect 5333 9216 5397 9220
rect 5413 9276 5477 9280
rect 5413 9220 5417 9276
rect 5417 9220 5473 9276
rect 5473 9220 5477 9276
rect 5413 9216 5477 9220
rect 5493 9276 5557 9280
rect 5493 9220 5497 9276
rect 5497 9220 5553 9276
rect 5553 9220 5557 9276
rect 5493 9216 5557 9220
rect 5573 9276 5637 9280
rect 5573 9220 5577 9276
rect 5577 9220 5633 9276
rect 5633 9220 5637 9276
rect 5573 9216 5637 9220
rect 8254 9276 8318 9280
rect 8254 9220 8258 9276
rect 8258 9220 8314 9276
rect 8314 9220 8318 9276
rect 8254 9216 8318 9220
rect 8334 9276 8398 9280
rect 8334 9220 8338 9276
rect 8338 9220 8394 9276
rect 8394 9220 8398 9276
rect 8334 9216 8398 9220
rect 8414 9276 8478 9280
rect 8414 9220 8418 9276
rect 8418 9220 8474 9276
rect 8474 9220 8478 9276
rect 8414 9216 8478 9220
rect 8494 9276 8558 9280
rect 8494 9220 8498 9276
rect 8498 9220 8554 9276
rect 8554 9220 8558 9276
rect 8494 9216 8558 9220
rect 11175 9276 11239 9280
rect 11175 9220 11179 9276
rect 11179 9220 11235 9276
rect 11235 9220 11239 9276
rect 11175 9216 11239 9220
rect 11255 9276 11319 9280
rect 11255 9220 11259 9276
rect 11259 9220 11315 9276
rect 11315 9220 11319 9276
rect 11255 9216 11319 9220
rect 11335 9276 11399 9280
rect 11335 9220 11339 9276
rect 11339 9220 11395 9276
rect 11395 9220 11399 9276
rect 11335 9216 11399 9220
rect 11415 9276 11479 9280
rect 11415 9220 11419 9276
rect 11419 9220 11475 9276
rect 11475 9220 11479 9276
rect 11415 9216 11479 9220
rect 3072 8732 3136 8736
rect 3072 8676 3076 8732
rect 3076 8676 3132 8732
rect 3132 8676 3136 8732
rect 3072 8672 3136 8676
rect 3152 8732 3216 8736
rect 3152 8676 3156 8732
rect 3156 8676 3212 8732
rect 3212 8676 3216 8732
rect 3152 8672 3216 8676
rect 3232 8732 3296 8736
rect 3232 8676 3236 8732
rect 3236 8676 3292 8732
rect 3292 8676 3296 8732
rect 3232 8672 3296 8676
rect 3312 8732 3376 8736
rect 3312 8676 3316 8732
rect 3316 8676 3372 8732
rect 3372 8676 3376 8732
rect 3312 8672 3376 8676
rect 5993 8732 6057 8736
rect 5993 8676 5997 8732
rect 5997 8676 6053 8732
rect 6053 8676 6057 8732
rect 5993 8672 6057 8676
rect 6073 8732 6137 8736
rect 6073 8676 6077 8732
rect 6077 8676 6133 8732
rect 6133 8676 6137 8732
rect 6073 8672 6137 8676
rect 6153 8732 6217 8736
rect 6153 8676 6157 8732
rect 6157 8676 6213 8732
rect 6213 8676 6217 8732
rect 6153 8672 6217 8676
rect 6233 8732 6297 8736
rect 6233 8676 6237 8732
rect 6237 8676 6293 8732
rect 6293 8676 6297 8732
rect 6233 8672 6297 8676
rect 8914 8732 8978 8736
rect 8914 8676 8918 8732
rect 8918 8676 8974 8732
rect 8974 8676 8978 8732
rect 8914 8672 8978 8676
rect 8994 8732 9058 8736
rect 8994 8676 8998 8732
rect 8998 8676 9054 8732
rect 9054 8676 9058 8732
rect 8994 8672 9058 8676
rect 9074 8732 9138 8736
rect 9074 8676 9078 8732
rect 9078 8676 9134 8732
rect 9134 8676 9138 8732
rect 9074 8672 9138 8676
rect 9154 8732 9218 8736
rect 9154 8676 9158 8732
rect 9158 8676 9214 8732
rect 9214 8676 9218 8732
rect 9154 8672 9218 8676
rect 11835 8732 11899 8736
rect 11835 8676 11839 8732
rect 11839 8676 11895 8732
rect 11895 8676 11899 8732
rect 11835 8672 11899 8676
rect 11915 8732 11979 8736
rect 11915 8676 11919 8732
rect 11919 8676 11975 8732
rect 11975 8676 11979 8732
rect 11915 8672 11979 8676
rect 11995 8732 12059 8736
rect 11995 8676 11999 8732
rect 11999 8676 12055 8732
rect 12055 8676 12059 8732
rect 11995 8672 12059 8676
rect 12075 8732 12139 8736
rect 12075 8676 12079 8732
rect 12079 8676 12135 8732
rect 12135 8676 12139 8732
rect 12075 8672 12139 8676
rect 2412 8188 2476 8192
rect 2412 8132 2416 8188
rect 2416 8132 2472 8188
rect 2472 8132 2476 8188
rect 2412 8128 2476 8132
rect 2492 8188 2556 8192
rect 2492 8132 2496 8188
rect 2496 8132 2552 8188
rect 2552 8132 2556 8188
rect 2492 8128 2556 8132
rect 2572 8188 2636 8192
rect 2572 8132 2576 8188
rect 2576 8132 2632 8188
rect 2632 8132 2636 8188
rect 2572 8128 2636 8132
rect 2652 8188 2716 8192
rect 2652 8132 2656 8188
rect 2656 8132 2712 8188
rect 2712 8132 2716 8188
rect 2652 8128 2716 8132
rect 5333 8188 5397 8192
rect 5333 8132 5337 8188
rect 5337 8132 5393 8188
rect 5393 8132 5397 8188
rect 5333 8128 5397 8132
rect 5413 8188 5477 8192
rect 5413 8132 5417 8188
rect 5417 8132 5473 8188
rect 5473 8132 5477 8188
rect 5413 8128 5477 8132
rect 5493 8188 5557 8192
rect 5493 8132 5497 8188
rect 5497 8132 5553 8188
rect 5553 8132 5557 8188
rect 5493 8128 5557 8132
rect 5573 8188 5637 8192
rect 5573 8132 5577 8188
rect 5577 8132 5633 8188
rect 5633 8132 5637 8188
rect 5573 8128 5637 8132
rect 8254 8188 8318 8192
rect 8254 8132 8258 8188
rect 8258 8132 8314 8188
rect 8314 8132 8318 8188
rect 8254 8128 8318 8132
rect 8334 8188 8398 8192
rect 8334 8132 8338 8188
rect 8338 8132 8394 8188
rect 8394 8132 8398 8188
rect 8334 8128 8398 8132
rect 8414 8188 8478 8192
rect 8414 8132 8418 8188
rect 8418 8132 8474 8188
rect 8474 8132 8478 8188
rect 8414 8128 8478 8132
rect 8494 8188 8558 8192
rect 8494 8132 8498 8188
rect 8498 8132 8554 8188
rect 8554 8132 8558 8188
rect 8494 8128 8558 8132
rect 11175 8188 11239 8192
rect 11175 8132 11179 8188
rect 11179 8132 11235 8188
rect 11235 8132 11239 8188
rect 11175 8128 11239 8132
rect 11255 8188 11319 8192
rect 11255 8132 11259 8188
rect 11259 8132 11315 8188
rect 11315 8132 11319 8188
rect 11255 8128 11319 8132
rect 11335 8188 11399 8192
rect 11335 8132 11339 8188
rect 11339 8132 11395 8188
rect 11395 8132 11399 8188
rect 11335 8128 11399 8132
rect 11415 8188 11479 8192
rect 11415 8132 11419 8188
rect 11419 8132 11475 8188
rect 11475 8132 11479 8188
rect 11415 8128 11479 8132
rect 3072 7644 3136 7648
rect 3072 7588 3076 7644
rect 3076 7588 3132 7644
rect 3132 7588 3136 7644
rect 3072 7584 3136 7588
rect 3152 7644 3216 7648
rect 3152 7588 3156 7644
rect 3156 7588 3212 7644
rect 3212 7588 3216 7644
rect 3152 7584 3216 7588
rect 3232 7644 3296 7648
rect 3232 7588 3236 7644
rect 3236 7588 3292 7644
rect 3292 7588 3296 7644
rect 3232 7584 3296 7588
rect 3312 7644 3376 7648
rect 3312 7588 3316 7644
rect 3316 7588 3372 7644
rect 3372 7588 3376 7644
rect 3312 7584 3376 7588
rect 5993 7644 6057 7648
rect 5993 7588 5997 7644
rect 5997 7588 6053 7644
rect 6053 7588 6057 7644
rect 5993 7584 6057 7588
rect 6073 7644 6137 7648
rect 6073 7588 6077 7644
rect 6077 7588 6133 7644
rect 6133 7588 6137 7644
rect 6073 7584 6137 7588
rect 6153 7644 6217 7648
rect 6153 7588 6157 7644
rect 6157 7588 6213 7644
rect 6213 7588 6217 7644
rect 6153 7584 6217 7588
rect 6233 7644 6297 7648
rect 6233 7588 6237 7644
rect 6237 7588 6293 7644
rect 6293 7588 6297 7644
rect 6233 7584 6297 7588
rect 8914 7644 8978 7648
rect 8914 7588 8918 7644
rect 8918 7588 8974 7644
rect 8974 7588 8978 7644
rect 8914 7584 8978 7588
rect 8994 7644 9058 7648
rect 8994 7588 8998 7644
rect 8998 7588 9054 7644
rect 9054 7588 9058 7644
rect 8994 7584 9058 7588
rect 9074 7644 9138 7648
rect 9074 7588 9078 7644
rect 9078 7588 9134 7644
rect 9134 7588 9138 7644
rect 9074 7584 9138 7588
rect 9154 7644 9218 7648
rect 9154 7588 9158 7644
rect 9158 7588 9214 7644
rect 9214 7588 9218 7644
rect 9154 7584 9218 7588
rect 11835 7644 11899 7648
rect 11835 7588 11839 7644
rect 11839 7588 11895 7644
rect 11895 7588 11899 7644
rect 11835 7584 11899 7588
rect 11915 7644 11979 7648
rect 11915 7588 11919 7644
rect 11919 7588 11975 7644
rect 11975 7588 11979 7644
rect 11915 7584 11979 7588
rect 11995 7644 12059 7648
rect 11995 7588 11999 7644
rect 11999 7588 12055 7644
rect 12055 7588 12059 7644
rect 11995 7584 12059 7588
rect 12075 7644 12139 7648
rect 12075 7588 12079 7644
rect 12079 7588 12135 7644
rect 12135 7588 12139 7644
rect 12075 7584 12139 7588
rect 2412 7100 2476 7104
rect 2412 7044 2416 7100
rect 2416 7044 2472 7100
rect 2472 7044 2476 7100
rect 2412 7040 2476 7044
rect 2492 7100 2556 7104
rect 2492 7044 2496 7100
rect 2496 7044 2552 7100
rect 2552 7044 2556 7100
rect 2492 7040 2556 7044
rect 2572 7100 2636 7104
rect 2572 7044 2576 7100
rect 2576 7044 2632 7100
rect 2632 7044 2636 7100
rect 2572 7040 2636 7044
rect 2652 7100 2716 7104
rect 2652 7044 2656 7100
rect 2656 7044 2712 7100
rect 2712 7044 2716 7100
rect 2652 7040 2716 7044
rect 5333 7100 5397 7104
rect 5333 7044 5337 7100
rect 5337 7044 5393 7100
rect 5393 7044 5397 7100
rect 5333 7040 5397 7044
rect 5413 7100 5477 7104
rect 5413 7044 5417 7100
rect 5417 7044 5473 7100
rect 5473 7044 5477 7100
rect 5413 7040 5477 7044
rect 5493 7100 5557 7104
rect 5493 7044 5497 7100
rect 5497 7044 5553 7100
rect 5553 7044 5557 7100
rect 5493 7040 5557 7044
rect 5573 7100 5637 7104
rect 5573 7044 5577 7100
rect 5577 7044 5633 7100
rect 5633 7044 5637 7100
rect 5573 7040 5637 7044
rect 8254 7100 8318 7104
rect 8254 7044 8258 7100
rect 8258 7044 8314 7100
rect 8314 7044 8318 7100
rect 8254 7040 8318 7044
rect 8334 7100 8398 7104
rect 8334 7044 8338 7100
rect 8338 7044 8394 7100
rect 8394 7044 8398 7100
rect 8334 7040 8398 7044
rect 8414 7100 8478 7104
rect 8414 7044 8418 7100
rect 8418 7044 8474 7100
rect 8474 7044 8478 7100
rect 8414 7040 8478 7044
rect 8494 7100 8558 7104
rect 8494 7044 8498 7100
rect 8498 7044 8554 7100
rect 8554 7044 8558 7100
rect 8494 7040 8558 7044
rect 11175 7100 11239 7104
rect 11175 7044 11179 7100
rect 11179 7044 11235 7100
rect 11235 7044 11239 7100
rect 11175 7040 11239 7044
rect 11255 7100 11319 7104
rect 11255 7044 11259 7100
rect 11259 7044 11315 7100
rect 11315 7044 11319 7100
rect 11255 7040 11319 7044
rect 11335 7100 11399 7104
rect 11335 7044 11339 7100
rect 11339 7044 11395 7100
rect 11395 7044 11399 7100
rect 11335 7040 11399 7044
rect 11415 7100 11479 7104
rect 11415 7044 11419 7100
rect 11419 7044 11475 7100
rect 11475 7044 11479 7100
rect 11415 7040 11479 7044
rect 3072 6556 3136 6560
rect 3072 6500 3076 6556
rect 3076 6500 3132 6556
rect 3132 6500 3136 6556
rect 3072 6496 3136 6500
rect 3152 6556 3216 6560
rect 3152 6500 3156 6556
rect 3156 6500 3212 6556
rect 3212 6500 3216 6556
rect 3152 6496 3216 6500
rect 3232 6556 3296 6560
rect 3232 6500 3236 6556
rect 3236 6500 3292 6556
rect 3292 6500 3296 6556
rect 3232 6496 3296 6500
rect 3312 6556 3376 6560
rect 3312 6500 3316 6556
rect 3316 6500 3372 6556
rect 3372 6500 3376 6556
rect 3312 6496 3376 6500
rect 5993 6556 6057 6560
rect 5993 6500 5997 6556
rect 5997 6500 6053 6556
rect 6053 6500 6057 6556
rect 5993 6496 6057 6500
rect 6073 6556 6137 6560
rect 6073 6500 6077 6556
rect 6077 6500 6133 6556
rect 6133 6500 6137 6556
rect 6073 6496 6137 6500
rect 6153 6556 6217 6560
rect 6153 6500 6157 6556
rect 6157 6500 6213 6556
rect 6213 6500 6217 6556
rect 6153 6496 6217 6500
rect 6233 6556 6297 6560
rect 6233 6500 6237 6556
rect 6237 6500 6293 6556
rect 6293 6500 6297 6556
rect 6233 6496 6297 6500
rect 8914 6556 8978 6560
rect 8914 6500 8918 6556
rect 8918 6500 8974 6556
rect 8974 6500 8978 6556
rect 8914 6496 8978 6500
rect 8994 6556 9058 6560
rect 8994 6500 8998 6556
rect 8998 6500 9054 6556
rect 9054 6500 9058 6556
rect 8994 6496 9058 6500
rect 9074 6556 9138 6560
rect 9074 6500 9078 6556
rect 9078 6500 9134 6556
rect 9134 6500 9138 6556
rect 9074 6496 9138 6500
rect 9154 6556 9218 6560
rect 9154 6500 9158 6556
rect 9158 6500 9214 6556
rect 9214 6500 9218 6556
rect 9154 6496 9218 6500
rect 11835 6556 11899 6560
rect 11835 6500 11839 6556
rect 11839 6500 11895 6556
rect 11895 6500 11899 6556
rect 11835 6496 11899 6500
rect 11915 6556 11979 6560
rect 11915 6500 11919 6556
rect 11919 6500 11975 6556
rect 11975 6500 11979 6556
rect 11915 6496 11979 6500
rect 11995 6556 12059 6560
rect 11995 6500 11999 6556
rect 11999 6500 12055 6556
rect 12055 6500 12059 6556
rect 11995 6496 12059 6500
rect 12075 6556 12139 6560
rect 12075 6500 12079 6556
rect 12079 6500 12135 6556
rect 12135 6500 12139 6556
rect 12075 6496 12139 6500
rect 2412 6012 2476 6016
rect 2412 5956 2416 6012
rect 2416 5956 2472 6012
rect 2472 5956 2476 6012
rect 2412 5952 2476 5956
rect 2492 6012 2556 6016
rect 2492 5956 2496 6012
rect 2496 5956 2552 6012
rect 2552 5956 2556 6012
rect 2492 5952 2556 5956
rect 2572 6012 2636 6016
rect 2572 5956 2576 6012
rect 2576 5956 2632 6012
rect 2632 5956 2636 6012
rect 2572 5952 2636 5956
rect 2652 6012 2716 6016
rect 2652 5956 2656 6012
rect 2656 5956 2712 6012
rect 2712 5956 2716 6012
rect 2652 5952 2716 5956
rect 5333 6012 5397 6016
rect 5333 5956 5337 6012
rect 5337 5956 5393 6012
rect 5393 5956 5397 6012
rect 5333 5952 5397 5956
rect 5413 6012 5477 6016
rect 5413 5956 5417 6012
rect 5417 5956 5473 6012
rect 5473 5956 5477 6012
rect 5413 5952 5477 5956
rect 5493 6012 5557 6016
rect 5493 5956 5497 6012
rect 5497 5956 5553 6012
rect 5553 5956 5557 6012
rect 5493 5952 5557 5956
rect 5573 6012 5637 6016
rect 5573 5956 5577 6012
rect 5577 5956 5633 6012
rect 5633 5956 5637 6012
rect 5573 5952 5637 5956
rect 8254 6012 8318 6016
rect 8254 5956 8258 6012
rect 8258 5956 8314 6012
rect 8314 5956 8318 6012
rect 8254 5952 8318 5956
rect 8334 6012 8398 6016
rect 8334 5956 8338 6012
rect 8338 5956 8394 6012
rect 8394 5956 8398 6012
rect 8334 5952 8398 5956
rect 8414 6012 8478 6016
rect 8414 5956 8418 6012
rect 8418 5956 8474 6012
rect 8474 5956 8478 6012
rect 8414 5952 8478 5956
rect 8494 6012 8558 6016
rect 8494 5956 8498 6012
rect 8498 5956 8554 6012
rect 8554 5956 8558 6012
rect 8494 5952 8558 5956
rect 11175 6012 11239 6016
rect 11175 5956 11179 6012
rect 11179 5956 11235 6012
rect 11235 5956 11239 6012
rect 11175 5952 11239 5956
rect 11255 6012 11319 6016
rect 11255 5956 11259 6012
rect 11259 5956 11315 6012
rect 11315 5956 11319 6012
rect 11255 5952 11319 5956
rect 11335 6012 11399 6016
rect 11335 5956 11339 6012
rect 11339 5956 11395 6012
rect 11395 5956 11399 6012
rect 11335 5952 11399 5956
rect 11415 6012 11479 6016
rect 11415 5956 11419 6012
rect 11419 5956 11475 6012
rect 11475 5956 11479 6012
rect 11415 5952 11479 5956
rect 3072 5468 3136 5472
rect 3072 5412 3076 5468
rect 3076 5412 3132 5468
rect 3132 5412 3136 5468
rect 3072 5408 3136 5412
rect 3152 5468 3216 5472
rect 3152 5412 3156 5468
rect 3156 5412 3212 5468
rect 3212 5412 3216 5468
rect 3152 5408 3216 5412
rect 3232 5468 3296 5472
rect 3232 5412 3236 5468
rect 3236 5412 3292 5468
rect 3292 5412 3296 5468
rect 3232 5408 3296 5412
rect 3312 5468 3376 5472
rect 3312 5412 3316 5468
rect 3316 5412 3372 5468
rect 3372 5412 3376 5468
rect 3312 5408 3376 5412
rect 5993 5468 6057 5472
rect 5993 5412 5997 5468
rect 5997 5412 6053 5468
rect 6053 5412 6057 5468
rect 5993 5408 6057 5412
rect 6073 5468 6137 5472
rect 6073 5412 6077 5468
rect 6077 5412 6133 5468
rect 6133 5412 6137 5468
rect 6073 5408 6137 5412
rect 6153 5468 6217 5472
rect 6153 5412 6157 5468
rect 6157 5412 6213 5468
rect 6213 5412 6217 5468
rect 6153 5408 6217 5412
rect 6233 5468 6297 5472
rect 6233 5412 6237 5468
rect 6237 5412 6293 5468
rect 6293 5412 6297 5468
rect 6233 5408 6297 5412
rect 8914 5468 8978 5472
rect 8914 5412 8918 5468
rect 8918 5412 8974 5468
rect 8974 5412 8978 5468
rect 8914 5408 8978 5412
rect 8994 5468 9058 5472
rect 8994 5412 8998 5468
rect 8998 5412 9054 5468
rect 9054 5412 9058 5468
rect 8994 5408 9058 5412
rect 9074 5468 9138 5472
rect 9074 5412 9078 5468
rect 9078 5412 9134 5468
rect 9134 5412 9138 5468
rect 9074 5408 9138 5412
rect 9154 5468 9218 5472
rect 9154 5412 9158 5468
rect 9158 5412 9214 5468
rect 9214 5412 9218 5468
rect 9154 5408 9218 5412
rect 11835 5468 11899 5472
rect 11835 5412 11839 5468
rect 11839 5412 11895 5468
rect 11895 5412 11899 5468
rect 11835 5408 11899 5412
rect 11915 5468 11979 5472
rect 11915 5412 11919 5468
rect 11919 5412 11975 5468
rect 11975 5412 11979 5468
rect 11915 5408 11979 5412
rect 11995 5468 12059 5472
rect 11995 5412 11999 5468
rect 11999 5412 12055 5468
rect 12055 5412 12059 5468
rect 11995 5408 12059 5412
rect 12075 5468 12139 5472
rect 12075 5412 12079 5468
rect 12079 5412 12135 5468
rect 12135 5412 12139 5468
rect 12075 5408 12139 5412
rect 2412 4924 2476 4928
rect 2412 4868 2416 4924
rect 2416 4868 2472 4924
rect 2472 4868 2476 4924
rect 2412 4864 2476 4868
rect 2492 4924 2556 4928
rect 2492 4868 2496 4924
rect 2496 4868 2552 4924
rect 2552 4868 2556 4924
rect 2492 4864 2556 4868
rect 2572 4924 2636 4928
rect 2572 4868 2576 4924
rect 2576 4868 2632 4924
rect 2632 4868 2636 4924
rect 2572 4864 2636 4868
rect 2652 4924 2716 4928
rect 2652 4868 2656 4924
rect 2656 4868 2712 4924
rect 2712 4868 2716 4924
rect 2652 4864 2716 4868
rect 5333 4924 5397 4928
rect 5333 4868 5337 4924
rect 5337 4868 5393 4924
rect 5393 4868 5397 4924
rect 5333 4864 5397 4868
rect 5413 4924 5477 4928
rect 5413 4868 5417 4924
rect 5417 4868 5473 4924
rect 5473 4868 5477 4924
rect 5413 4864 5477 4868
rect 5493 4924 5557 4928
rect 5493 4868 5497 4924
rect 5497 4868 5553 4924
rect 5553 4868 5557 4924
rect 5493 4864 5557 4868
rect 5573 4924 5637 4928
rect 5573 4868 5577 4924
rect 5577 4868 5633 4924
rect 5633 4868 5637 4924
rect 5573 4864 5637 4868
rect 8254 4924 8318 4928
rect 8254 4868 8258 4924
rect 8258 4868 8314 4924
rect 8314 4868 8318 4924
rect 8254 4864 8318 4868
rect 8334 4924 8398 4928
rect 8334 4868 8338 4924
rect 8338 4868 8394 4924
rect 8394 4868 8398 4924
rect 8334 4864 8398 4868
rect 8414 4924 8478 4928
rect 8414 4868 8418 4924
rect 8418 4868 8474 4924
rect 8474 4868 8478 4924
rect 8414 4864 8478 4868
rect 8494 4924 8558 4928
rect 8494 4868 8498 4924
rect 8498 4868 8554 4924
rect 8554 4868 8558 4924
rect 8494 4864 8558 4868
rect 11175 4924 11239 4928
rect 11175 4868 11179 4924
rect 11179 4868 11235 4924
rect 11235 4868 11239 4924
rect 11175 4864 11239 4868
rect 11255 4924 11319 4928
rect 11255 4868 11259 4924
rect 11259 4868 11315 4924
rect 11315 4868 11319 4924
rect 11255 4864 11319 4868
rect 11335 4924 11399 4928
rect 11335 4868 11339 4924
rect 11339 4868 11395 4924
rect 11395 4868 11399 4924
rect 11335 4864 11399 4868
rect 11415 4924 11479 4928
rect 11415 4868 11419 4924
rect 11419 4868 11475 4924
rect 11475 4868 11479 4924
rect 11415 4864 11479 4868
rect 3072 4380 3136 4384
rect 3072 4324 3076 4380
rect 3076 4324 3132 4380
rect 3132 4324 3136 4380
rect 3072 4320 3136 4324
rect 3152 4380 3216 4384
rect 3152 4324 3156 4380
rect 3156 4324 3212 4380
rect 3212 4324 3216 4380
rect 3152 4320 3216 4324
rect 3232 4380 3296 4384
rect 3232 4324 3236 4380
rect 3236 4324 3292 4380
rect 3292 4324 3296 4380
rect 3232 4320 3296 4324
rect 3312 4380 3376 4384
rect 3312 4324 3316 4380
rect 3316 4324 3372 4380
rect 3372 4324 3376 4380
rect 3312 4320 3376 4324
rect 5993 4380 6057 4384
rect 5993 4324 5997 4380
rect 5997 4324 6053 4380
rect 6053 4324 6057 4380
rect 5993 4320 6057 4324
rect 6073 4380 6137 4384
rect 6073 4324 6077 4380
rect 6077 4324 6133 4380
rect 6133 4324 6137 4380
rect 6073 4320 6137 4324
rect 6153 4380 6217 4384
rect 6153 4324 6157 4380
rect 6157 4324 6213 4380
rect 6213 4324 6217 4380
rect 6153 4320 6217 4324
rect 6233 4380 6297 4384
rect 6233 4324 6237 4380
rect 6237 4324 6293 4380
rect 6293 4324 6297 4380
rect 6233 4320 6297 4324
rect 8914 4380 8978 4384
rect 8914 4324 8918 4380
rect 8918 4324 8974 4380
rect 8974 4324 8978 4380
rect 8914 4320 8978 4324
rect 8994 4380 9058 4384
rect 8994 4324 8998 4380
rect 8998 4324 9054 4380
rect 9054 4324 9058 4380
rect 8994 4320 9058 4324
rect 9074 4380 9138 4384
rect 9074 4324 9078 4380
rect 9078 4324 9134 4380
rect 9134 4324 9138 4380
rect 9074 4320 9138 4324
rect 9154 4380 9218 4384
rect 9154 4324 9158 4380
rect 9158 4324 9214 4380
rect 9214 4324 9218 4380
rect 9154 4320 9218 4324
rect 11835 4380 11899 4384
rect 11835 4324 11839 4380
rect 11839 4324 11895 4380
rect 11895 4324 11899 4380
rect 11835 4320 11899 4324
rect 11915 4380 11979 4384
rect 11915 4324 11919 4380
rect 11919 4324 11975 4380
rect 11975 4324 11979 4380
rect 11915 4320 11979 4324
rect 11995 4380 12059 4384
rect 11995 4324 11999 4380
rect 11999 4324 12055 4380
rect 12055 4324 12059 4380
rect 11995 4320 12059 4324
rect 12075 4380 12139 4384
rect 12075 4324 12079 4380
rect 12079 4324 12135 4380
rect 12135 4324 12139 4380
rect 12075 4320 12139 4324
rect 2412 3836 2476 3840
rect 2412 3780 2416 3836
rect 2416 3780 2472 3836
rect 2472 3780 2476 3836
rect 2412 3776 2476 3780
rect 2492 3836 2556 3840
rect 2492 3780 2496 3836
rect 2496 3780 2552 3836
rect 2552 3780 2556 3836
rect 2492 3776 2556 3780
rect 2572 3836 2636 3840
rect 2572 3780 2576 3836
rect 2576 3780 2632 3836
rect 2632 3780 2636 3836
rect 2572 3776 2636 3780
rect 2652 3836 2716 3840
rect 2652 3780 2656 3836
rect 2656 3780 2712 3836
rect 2712 3780 2716 3836
rect 2652 3776 2716 3780
rect 5333 3836 5397 3840
rect 5333 3780 5337 3836
rect 5337 3780 5393 3836
rect 5393 3780 5397 3836
rect 5333 3776 5397 3780
rect 5413 3836 5477 3840
rect 5413 3780 5417 3836
rect 5417 3780 5473 3836
rect 5473 3780 5477 3836
rect 5413 3776 5477 3780
rect 5493 3836 5557 3840
rect 5493 3780 5497 3836
rect 5497 3780 5553 3836
rect 5553 3780 5557 3836
rect 5493 3776 5557 3780
rect 5573 3836 5637 3840
rect 5573 3780 5577 3836
rect 5577 3780 5633 3836
rect 5633 3780 5637 3836
rect 5573 3776 5637 3780
rect 8254 3836 8318 3840
rect 8254 3780 8258 3836
rect 8258 3780 8314 3836
rect 8314 3780 8318 3836
rect 8254 3776 8318 3780
rect 8334 3836 8398 3840
rect 8334 3780 8338 3836
rect 8338 3780 8394 3836
rect 8394 3780 8398 3836
rect 8334 3776 8398 3780
rect 8414 3836 8478 3840
rect 8414 3780 8418 3836
rect 8418 3780 8474 3836
rect 8474 3780 8478 3836
rect 8414 3776 8478 3780
rect 8494 3836 8558 3840
rect 8494 3780 8498 3836
rect 8498 3780 8554 3836
rect 8554 3780 8558 3836
rect 8494 3776 8558 3780
rect 11175 3836 11239 3840
rect 11175 3780 11179 3836
rect 11179 3780 11235 3836
rect 11235 3780 11239 3836
rect 11175 3776 11239 3780
rect 11255 3836 11319 3840
rect 11255 3780 11259 3836
rect 11259 3780 11315 3836
rect 11315 3780 11319 3836
rect 11255 3776 11319 3780
rect 11335 3836 11399 3840
rect 11335 3780 11339 3836
rect 11339 3780 11395 3836
rect 11395 3780 11399 3836
rect 11335 3776 11399 3780
rect 11415 3836 11479 3840
rect 11415 3780 11419 3836
rect 11419 3780 11475 3836
rect 11475 3780 11479 3836
rect 11415 3776 11479 3780
rect 3072 3292 3136 3296
rect 3072 3236 3076 3292
rect 3076 3236 3132 3292
rect 3132 3236 3136 3292
rect 3072 3232 3136 3236
rect 3152 3292 3216 3296
rect 3152 3236 3156 3292
rect 3156 3236 3212 3292
rect 3212 3236 3216 3292
rect 3152 3232 3216 3236
rect 3232 3292 3296 3296
rect 3232 3236 3236 3292
rect 3236 3236 3292 3292
rect 3292 3236 3296 3292
rect 3232 3232 3296 3236
rect 3312 3292 3376 3296
rect 3312 3236 3316 3292
rect 3316 3236 3372 3292
rect 3372 3236 3376 3292
rect 3312 3232 3376 3236
rect 5993 3292 6057 3296
rect 5993 3236 5997 3292
rect 5997 3236 6053 3292
rect 6053 3236 6057 3292
rect 5993 3232 6057 3236
rect 6073 3292 6137 3296
rect 6073 3236 6077 3292
rect 6077 3236 6133 3292
rect 6133 3236 6137 3292
rect 6073 3232 6137 3236
rect 6153 3292 6217 3296
rect 6153 3236 6157 3292
rect 6157 3236 6213 3292
rect 6213 3236 6217 3292
rect 6153 3232 6217 3236
rect 6233 3292 6297 3296
rect 6233 3236 6237 3292
rect 6237 3236 6293 3292
rect 6293 3236 6297 3292
rect 6233 3232 6297 3236
rect 8914 3292 8978 3296
rect 8914 3236 8918 3292
rect 8918 3236 8974 3292
rect 8974 3236 8978 3292
rect 8914 3232 8978 3236
rect 8994 3292 9058 3296
rect 8994 3236 8998 3292
rect 8998 3236 9054 3292
rect 9054 3236 9058 3292
rect 8994 3232 9058 3236
rect 9074 3292 9138 3296
rect 9074 3236 9078 3292
rect 9078 3236 9134 3292
rect 9134 3236 9138 3292
rect 9074 3232 9138 3236
rect 9154 3292 9218 3296
rect 9154 3236 9158 3292
rect 9158 3236 9214 3292
rect 9214 3236 9218 3292
rect 9154 3232 9218 3236
rect 11835 3292 11899 3296
rect 11835 3236 11839 3292
rect 11839 3236 11895 3292
rect 11895 3236 11899 3292
rect 11835 3232 11899 3236
rect 11915 3292 11979 3296
rect 11915 3236 11919 3292
rect 11919 3236 11975 3292
rect 11975 3236 11979 3292
rect 11915 3232 11979 3236
rect 11995 3292 12059 3296
rect 11995 3236 11999 3292
rect 11999 3236 12055 3292
rect 12055 3236 12059 3292
rect 11995 3232 12059 3236
rect 12075 3292 12139 3296
rect 12075 3236 12079 3292
rect 12079 3236 12135 3292
rect 12135 3236 12139 3292
rect 12075 3232 12139 3236
rect 2412 2748 2476 2752
rect 2412 2692 2416 2748
rect 2416 2692 2472 2748
rect 2472 2692 2476 2748
rect 2412 2688 2476 2692
rect 2492 2748 2556 2752
rect 2492 2692 2496 2748
rect 2496 2692 2552 2748
rect 2552 2692 2556 2748
rect 2492 2688 2556 2692
rect 2572 2748 2636 2752
rect 2572 2692 2576 2748
rect 2576 2692 2632 2748
rect 2632 2692 2636 2748
rect 2572 2688 2636 2692
rect 2652 2748 2716 2752
rect 2652 2692 2656 2748
rect 2656 2692 2712 2748
rect 2712 2692 2716 2748
rect 2652 2688 2716 2692
rect 5333 2748 5397 2752
rect 5333 2692 5337 2748
rect 5337 2692 5393 2748
rect 5393 2692 5397 2748
rect 5333 2688 5397 2692
rect 5413 2748 5477 2752
rect 5413 2692 5417 2748
rect 5417 2692 5473 2748
rect 5473 2692 5477 2748
rect 5413 2688 5477 2692
rect 5493 2748 5557 2752
rect 5493 2692 5497 2748
rect 5497 2692 5553 2748
rect 5553 2692 5557 2748
rect 5493 2688 5557 2692
rect 5573 2748 5637 2752
rect 5573 2692 5577 2748
rect 5577 2692 5633 2748
rect 5633 2692 5637 2748
rect 5573 2688 5637 2692
rect 8254 2748 8318 2752
rect 8254 2692 8258 2748
rect 8258 2692 8314 2748
rect 8314 2692 8318 2748
rect 8254 2688 8318 2692
rect 8334 2748 8398 2752
rect 8334 2692 8338 2748
rect 8338 2692 8394 2748
rect 8394 2692 8398 2748
rect 8334 2688 8398 2692
rect 8414 2748 8478 2752
rect 8414 2692 8418 2748
rect 8418 2692 8474 2748
rect 8474 2692 8478 2748
rect 8414 2688 8478 2692
rect 8494 2748 8558 2752
rect 8494 2692 8498 2748
rect 8498 2692 8554 2748
rect 8554 2692 8558 2748
rect 8494 2688 8558 2692
rect 11175 2748 11239 2752
rect 11175 2692 11179 2748
rect 11179 2692 11235 2748
rect 11235 2692 11239 2748
rect 11175 2688 11239 2692
rect 11255 2748 11319 2752
rect 11255 2692 11259 2748
rect 11259 2692 11315 2748
rect 11315 2692 11319 2748
rect 11255 2688 11319 2692
rect 11335 2748 11399 2752
rect 11335 2692 11339 2748
rect 11339 2692 11395 2748
rect 11395 2692 11399 2748
rect 11335 2688 11399 2692
rect 11415 2748 11479 2752
rect 11415 2692 11419 2748
rect 11419 2692 11475 2748
rect 11475 2692 11479 2748
rect 11415 2688 11479 2692
rect 3072 2204 3136 2208
rect 3072 2148 3076 2204
rect 3076 2148 3132 2204
rect 3132 2148 3136 2204
rect 3072 2144 3136 2148
rect 3152 2204 3216 2208
rect 3152 2148 3156 2204
rect 3156 2148 3212 2204
rect 3212 2148 3216 2204
rect 3152 2144 3216 2148
rect 3232 2204 3296 2208
rect 3232 2148 3236 2204
rect 3236 2148 3292 2204
rect 3292 2148 3296 2204
rect 3232 2144 3296 2148
rect 3312 2204 3376 2208
rect 3312 2148 3316 2204
rect 3316 2148 3372 2204
rect 3372 2148 3376 2204
rect 3312 2144 3376 2148
rect 5993 2204 6057 2208
rect 5993 2148 5997 2204
rect 5997 2148 6053 2204
rect 6053 2148 6057 2204
rect 5993 2144 6057 2148
rect 6073 2204 6137 2208
rect 6073 2148 6077 2204
rect 6077 2148 6133 2204
rect 6133 2148 6137 2204
rect 6073 2144 6137 2148
rect 6153 2204 6217 2208
rect 6153 2148 6157 2204
rect 6157 2148 6213 2204
rect 6213 2148 6217 2204
rect 6153 2144 6217 2148
rect 6233 2204 6297 2208
rect 6233 2148 6237 2204
rect 6237 2148 6293 2204
rect 6293 2148 6297 2204
rect 6233 2144 6297 2148
rect 8914 2204 8978 2208
rect 8914 2148 8918 2204
rect 8918 2148 8974 2204
rect 8974 2148 8978 2204
rect 8914 2144 8978 2148
rect 8994 2204 9058 2208
rect 8994 2148 8998 2204
rect 8998 2148 9054 2204
rect 9054 2148 9058 2204
rect 8994 2144 9058 2148
rect 9074 2204 9138 2208
rect 9074 2148 9078 2204
rect 9078 2148 9134 2204
rect 9134 2148 9138 2204
rect 9074 2144 9138 2148
rect 9154 2204 9218 2208
rect 9154 2148 9158 2204
rect 9158 2148 9214 2204
rect 9214 2148 9218 2204
rect 9154 2144 9218 2148
rect 11835 2204 11899 2208
rect 11835 2148 11839 2204
rect 11839 2148 11895 2204
rect 11895 2148 11899 2204
rect 11835 2144 11899 2148
rect 11915 2204 11979 2208
rect 11915 2148 11919 2204
rect 11919 2148 11975 2204
rect 11975 2148 11979 2204
rect 11915 2144 11979 2148
rect 11995 2204 12059 2208
rect 11995 2148 11999 2204
rect 11999 2148 12055 2204
rect 12055 2148 12059 2204
rect 11995 2144 12059 2148
rect 12075 2204 12139 2208
rect 12075 2148 12079 2204
rect 12079 2148 12135 2204
rect 12135 2148 12139 2204
rect 12075 2144 12139 2148
<< metal4 >>
rect 2404 13632 2724 13648
rect 2404 13568 2412 13632
rect 2476 13568 2492 13632
rect 2556 13568 2572 13632
rect 2636 13568 2652 13632
rect 2716 13568 2724 13632
rect 2404 12544 2724 13568
rect 2404 12480 2412 12544
rect 2476 12480 2492 12544
rect 2556 12480 2572 12544
rect 2636 12480 2652 12544
rect 2716 12480 2724 12544
rect 2404 12290 2724 12480
rect 2404 12054 2446 12290
rect 2682 12054 2724 12290
rect 2404 11456 2724 12054
rect 2404 11392 2412 11456
rect 2476 11392 2492 11456
rect 2556 11392 2572 11456
rect 2636 11392 2652 11456
rect 2716 11392 2724 11456
rect 2404 10368 2724 11392
rect 2404 10304 2412 10368
rect 2476 10304 2492 10368
rect 2556 10304 2572 10368
rect 2636 10304 2652 10368
rect 2716 10304 2724 10368
rect 2404 9434 2724 10304
rect 2404 9280 2446 9434
rect 2682 9280 2724 9434
rect 2404 9216 2412 9280
rect 2716 9216 2724 9280
rect 2404 9198 2446 9216
rect 2682 9198 2724 9216
rect 2404 8192 2724 9198
rect 2404 8128 2412 8192
rect 2476 8128 2492 8192
rect 2556 8128 2572 8192
rect 2636 8128 2652 8192
rect 2716 8128 2724 8192
rect 2404 7104 2724 8128
rect 2404 7040 2412 7104
rect 2476 7040 2492 7104
rect 2556 7040 2572 7104
rect 2636 7040 2652 7104
rect 2716 7040 2724 7104
rect 2404 6578 2724 7040
rect 2404 6342 2446 6578
rect 2682 6342 2724 6578
rect 2404 6016 2724 6342
rect 2404 5952 2412 6016
rect 2476 5952 2492 6016
rect 2556 5952 2572 6016
rect 2636 5952 2652 6016
rect 2716 5952 2724 6016
rect 2404 4928 2724 5952
rect 2404 4864 2412 4928
rect 2476 4864 2492 4928
rect 2556 4864 2572 4928
rect 2636 4864 2652 4928
rect 2716 4864 2724 4928
rect 2404 3840 2724 4864
rect 2404 3776 2412 3840
rect 2476 3776 2492 3840
rect 2556 3776 2572 3840
rect 2636 3776 2652 3840
rect 2716 3776 2724 3840
rect 2404 3722 2724 3776
rect 2404 3486 2446 3722
rect 2682 3486 2724 3722
rect 2404 2752 2724 3486
rect 2404 2688 2412 2752
rect 2476 2688 2492 2752
rect 2556 2688 2572 2752
rect 2636 2688 2652 2752
rect 2716 2688 2724 2752
rect 2404 2128 2724 2688
rect 3064 13088 3384 13648
rect 3064 13024 3072 13088
rect 3136 13024 3152 13088
rect 3216 13024 3232 13088
rect 3296 13024 3312 13088
rect 3376 13024 3384 13088
rect 3064 12950 3384 13024
rect 3064 12714 3106 12950
rect 3342 12714 3384 12950
rect 3064 12000 3384 12714
rect 3064 11936 3072 12000
rect 3136 11936 3152 12000
rect 3216 11936 3232 12000
rect 3296 11936 3312 12000
rect 3376 11936 3384 12000
rect 3064 10912 3384 11936
rect 3064 10848 3072 10912
rect 3136 10848 3152 10912
rect 3216 10848 3232 10912
rect 3296 10848 3312 10912
rect 3376 10848 3384 10912
rect 3064 10094 3384 10848
rect 3064 9858 3106 10094
rect 3342 9858 3384 10094
rect 3064 9824 3384 9858
rect 3064 9760 3072 9824
rect 3136 9760 3152 9824
rect 3216 9760 3232 9824
rect 3296 9760 3312 9824
rect 3376 9760 3384 9824
rect 3064 8736 3384 9760
rect 3064 8672 3072 8736
rect 3136 8672 3152 8736
rect 3216 8672 3232 8736
rect 3296 8672 3312 8736
rect 3376 8672 3384 8736
rect 3064 7648 3384 8672
rect 3064 7584 3072 7648
rect 3136 7584 3152 7648
rect 3216 7584 3232 7648
rect 3296 7584 3312 7648
rect 3376 7584 3384 7648
rect 3064 7238 3384 7584
rect 3064 7002 3106 7238
rect 3342 7002 3384 7238
rect 3064 6560 3384 7002
rect 3064 6496 3072 6560
rect 3136 6496 3152 6560
rect 3216 6496 3232 6560
rect 3296 6496 3312 6560
rect 3376 6496 3384 6560
rect 3064 5472 3384 6496
rect 3064 5408 3072 5472
rect 3136 5408 3152 5472
rect 3216 5408 3232 5472
rect 3296 5408 3312 5472
rect 3376 5408 3384 5472
rect 3064 4384 3384 5408
rect 3064 4320 3072 4384
rect 3136 4382 3152 4384
rect 3216 4382 3232 4384
rect 3296 4382 3312 4384
rect 3376 4320 3384 4384
rect 3064 4146 3106 4320
rect 3342 4146 3384 4320
rect 3064 3296 3384 4146
rect 3064 3232 3072 3296
rect 3136 3232 3152 3296
rect 3216 3232 3232 3296
rect 3296 3232 3312 3296
rect 3376 3232 3384 3296
rect 3064 2208 3384 3232
rect 3064 2144 3072 2208
rect 3136 2144 3152 2208
rect 3216 2144 3232 2208
rect 3296 2144 3312 2208
rect 3376 2144 3384 2208
rect 3064 2128 3384 2144
rect 5325 13632 5645 13648
rect 5325 13568 5333 13632
rect 5397 13568 5413 13632
rect 5477 13568 5493 13632
rect 5557 13568 5573 13632
rect 5637 13568 5645 13632
rect 5325 12544 5645 13568
rect 5325 12480 5333 12544
rect 5397 12480 5413 12544
rect 5477 12480 5493 12544
rect 5557 12480 5573 12544
rect 5637 12480 5645 12544
rect 5325 12290 5645 12480
rect 5325 12054 5367 12290
rect 5603 12054 5645 12290
rect 5325 11456 5645 12054
rect 5325 11392 5333 11456
rect 5397 11392 5413 11456
rect 5477 11392 5493 11456
rect 5557 11392 5573 11456
rect 5637 11392 5645 11456
rect 5325 10368 5645 11392
rect 5325 10304 5333 10368
rect 5397 10304 5413 10368
rect 5477 10304 5493 10368
rect 5557 10304 5573 10368
rect 5637 10304 5645 10368
rect 5325 9434 5645 10304
rect 5325 9280 5367 9434
rect 5603 9280 5645 9434
rect 5325 9216 5333 9280
rect 5637 9216 5645 9280
rect 5325 9198 5367 9216
rect 5603 9198 5645 9216
rect 5325 8192 5645 9198
rect 5325 8128 5333 8192
rect 5397 8128 5413 8192
rect 5477 8128 5493 8192
rect 5557 8128 5573 8192
rect 5637 8128 5645 8192
rect 5325 7104 5645 8128
rect 5325 7040 5333 7104
rect 5397 7040 5413 7104
rect 5477 7040 5493 7104
rect 5557 7040 5573 7104
rect 5637 7040 5645 7104
rect 5325 6578 5645 7040
rect 5325 6342 5367 6578
rect 5603 6342 5645 6578
rect 5325 6016 5645 6342
rect 5325 5952 5333 6016
rect 5397 5952 5413 6016
rect 5477 5952 5493 6016
rect 5557 5952 5573 6016
rect 5637 5952 5645 6016
rect 5325 4928 5645 5952
rect 5325 4864 5333 4928
rect 5397 4864 5413 4928
rect 5477 4864 5493 4928
rect 5557 4864 5573 4928
rect 5637 4864 5645 4928
rect 5325 3840 5645 4864
rect 5325 3776 5333 3840
rect 5397 3776 5413 3840
rect 5477 3776 5493 3840
rect 5557 3776 5573 3840
rect 5637 3776 5645 3840
rect 5325 3722 5645 3776
rect 5325 3486 5367 3722
rect 5603 3486 5645 3722
rect 5325 2752 5645 3486
rect 5325 2688 5333 2752
rect 5397 2688 5413 2752
rect 5477 2688 5493 2752
rect 5557 2688 5573 2752
rect 5637 2688 5645 2752
rect 5325 2128 5645 2688
rect 5985 13088 6305 13648
rect 5985 13024 5993 13088
rect 6057 13024 6073 13088
rect 6137 13024 6153 13088
rect 6217 13024 6233 13088
rect 6297 13024 6305 13088
rect 5985 12950 6305 13024
rect 5985 12714 6027 12950
rect 6263 12714 6305 12950
rect 5985 12000 6305 12714
rect 5985 11936 5993 12000
rect 6057 11936 6073 12000
rect 6137 11936 6153 12000
rect 6217 11936 6233 12000
rect 6297 11936 6305 12000
rect 5985 10912 6305 11936
rect 5985 10848 5993 10912
rect 6057 10848 6073 10912
rect 6137 10848 6153 10912
rect 6217 10848 6233 10912
rect 6297 10848 6305 10912
rect 5985 10094 6305 10848
rect 5985 9858 6027 10094
rect 6263 9858 6305 10094
rect 5985 9824 6305 9858
rect 5985 9760 5993 9824
rect 6057 9760 6073 9824
rect 6137 9760 6153 9824
rect 6217 9760 6233 9824
rect 6297 9760 6305 9824
rect 5985 8736 6305 9760
rect 5985 8672 5993 8736
rect 6057 8672 6073 8736
rect 6137 8672 6153 8736
rect 6217 8672 6233 8736
rect 6297 8672 6305 8736
rect 5985 7648 6305 8672
rect 5985 7584 5993 7648
rect 6057 7584 6073 7648
rect 6137 7584 6153 7648
rect 6217 7584 6233 7648
rect 6297 7584 6305 7648
rect 5985 7238 6305 7584
rect 5985 7002 6027 7238
rect 6263 7002 6305 7238
rect 5985 6560 6305 7002
rect 5985 6496 5993 6560
rect 6057 6496 6073 6560
rect 6137 6496 6153 6560
rect 6217 6496 6233 6560
rect 6297 6496 6305 6560
rect 5985 5472 6305 6496
rect 5985 5408 5993 5472
rect 6057 5408 6073 5472
rect 6137 5408 6153 5472
rect 6217 5408 6233 5472
rect 6297 5408 6305 5472
rect 5985 4384 6305 5408
rect 5985 4320 5993 4384
rect 6057 4382 6073 4384
rect 6137 4382 6153 4384
rect 6217 4382 6233 4384
rect 6297 4320 6305 4384
rect 5985 4146 6027 4320
rect 6263 4146 6305 4320
rect 5985 3296 6305 4146
rect 5985 3232 5993 3296
rect 6057 3232 6073 3296
rect 6137 3232 6153 3296
rect 6217 3232 6233 3296
rect 6297 3232 6305 3296
rect 5985 2208 6305 3232
rect 5985 2144 5993 2208
rect 6057 2144 6073 2208
rect 6137 2144 6153 2208
rect 6217 2144 6233 2208
rect 6297 2144 6305 2208
rect 5985 2128 6305 2144
rect 8246 13632 8566 13648
rect 8246 13568 8254 13632
rect 8318 13568 8334 13632
rect 8398 13568 8414 13632
rect 8478 13568 8494 13632
rect 8558 13568 8566 13632
rect 8246 12544 8566 13568
rect 8246 12480 8254 12544
rect 8318 12480 8334 12544
rect 8398 12480 8414 12544
rect 8478 12480 8494 12544
rect 8558 12480 8566 12544
rect 8246 12290 8566 12480
rect 8246 12054 8288 12290
rect 8524 12054 8566 12290
rect 8246 11456 8566 12054
rect 8246 11392 8254 11456
rect 8318 11392 8334 11456
rect 8398 11392 8414 11456
rect 8478 11392 8494 11456
rect 8558 11392 8566 11456
rect 8246 10368 8566 11392
rect 8246 10304 8254 10368
rect 8318 10304 8334 10368
rect 8398 10304 8414 10368
rect 8478 10304 8494 10368
rect 8558 10304 8566 10368
rect 8246 9434 8566 10304
rect 8246 9280 8288 9434
rect 8524 9280 8566 9434
rect 8246 9216 8254 9280
rect 8558 9216 8566 9280
rect 8246 9198 8288 9216
rect 8524 9198 8566 9216
rect 8246 8192 8566 9198
rect 8246 8128 8254 8192
rect 8318 8128 8334 8192
rect 8398 8128 8414 8192
rect 8478 8128 8494 8192
rect 8558 8128 8566 8192
rect 8246 7104 8566 8128
rect 8246 7040 8254 7104
rect 8318 7040 8334 7104
rect 8398 7040 8414 7104
rect 8478 7040 8494 7104
rect 8558 7040 8566 7104
rect 8246 6578 8566 7040
rect 8246 6342 8288 6578
rect 8524 6342 8566 6578
rect 8246 6016 8566 6342
rect 8246 5952 8254 6016
rect 8318 5952 8334 6016
rect 8398 5952 8414 6016
rect 8478 5952 8494 6016
rect 8558 5952 8566 6016
rect 8246 4928 8566 5952
rect 8246 4864 8254 4928
rect 8318 4864 8334 4928
rect 8398 4864 8414 4928
rect 8478 4864 8494 4928
rect 8558 4864 8566 4928
rect 8246 3840 8566 4864
rect 8246 3776 8254 3840
rect 8318 3776 8334 3840
rect 8398 3776 8414 3840
rect 8478 3776 8494 3840
rect 8558 3776 8566 3840
rect 8246 3722 8566 3776
rect 8246 3486 8288 3722
rect 8524 3486 8566 3722
rect 8246 2752 8566 3486
rect 8246 2688 8254 2752
rect 8318 2688 8334 2752
rect 8398 2688 8414 2752
rect 8478 2688 8494 2752
rect 8558 2688 8566 2752
rect 8246 2128 8566 2688
rect 8906 13088 9226 13648
rect 8906 13024 8914 13088
rect 8978 13024 8994 13088
rect 9058 13024 9074 13088
rect 9138 13024 9154 13088
rect 9218 13024 9226 13088
rect 8906 12950 9226 13024
rect 8906 12714 8948 12950
rect 9184 12714 9226 12950
rect 8906 12000 9226 12714
rect 8906 11936 8914 12000
rect 8978 11936 8994 12000
rect 9058 11936 9074 12000
rect 9138 11936 9154 12000
rect 9218 11936 9226 12000
rect 8906 10912 9226 11936
rect 8906 10848 8914 10912
rect 8978 10848 8994 10912
rect 9058 10848 9074 10912
rect 9138 10848 9154 10912
rect 9218 10848 9226 10912
rect 8906 10094 9226 10848
rect 8906 9858 8948 10094
rect 9184 9858 9226 10094
rect 8906 9824 9226 9858
rect 8906 9760 8914 9824
rect 8978 9760 8994 9824
rect 9058 9760 9074 9824
rect 9138 9760 9154 9824
rect 9218 9760 9226 9824
rect 8906 8736 9226 9760
rect 8906 8672 8914 8736
rect 8978 8672 8994 8736
rect 9058 8672 9074 8736
rect 9138 8672 9154 8736
rect 9218 8672 9226 8736
rect 8906 7648 9226 8672
rect 8906 7584 8914 7648
rect 8978 7584 8994 7648
rect 9058 7584 9074 7648
rect 9138 7584 9154 7648
rect 9218 7584 9226 7648
rect 8906 7238 9226 7584
rect 8906 7002 8948 7238
rect 9184 7002 9226 7238
rect 8906 6560 9226 7002
rect 8906 6496 8914 6560
rect 8978 6496 8994 6560
rect 9058 6496 9074 6560
rect 9138 6496 9154 6560
rect 9218 6496 9226 6560
rect 8906 5472 9226 6496
rect 8906 5408 8914 5472
rect 8978 5408 8994 5472
rect 9058 5408 9074 5472
rect 9138 5408 9154 5472
rect 9218 5408 9226 5472
rect 8906 4384 9226 5408
rect 8906 4320 8914 4384
rect 8978 4382 8994 4384
rect 9058 4382 9074 4384
rect 9138 4382 9154 4384
rect 9218 4320 9226 4384
rect 8906 4146 8948 4320
rect 9184 4146 9226 4320
rect 8906 3296 9226 4146
rect 8906 3232 8914 3296
rect 8978 3232 8994 3296
rect 9058 3232 9074 3296
rect 9138 3232 9154 3296
rect 9218 3232 9226 3296
rect 8906 2208 9226 3232
rect 8906 2144 8914 2208
rect 8978 2144 8994 2208
rect 9058 2144 9074 2208
rect 9138 2144 9154 2208
rect 9218 2144 9226 2208
rect 8906 2128 9226 2144
rect 11167 13632 11487 13648
rect 11167 13568 11175 13632
rect 11239 13568 11255 13632
rect 11319 13568 11335 13632
rect 11399 13568 11415 13632
rect 11479 13568 11487 13632
rect 11167 12544 11487 13568
rect 11167 12480 11175 12544
rect 11239 12480 11255 12544
rect 11319 12480 11335 12544
rect 11399 12480 11415 12544
rect 11479 12480 11487 12544
rect 11167 12290 11487 12480
rect 11167 12054 11209 12290
rect 11445 12054 11487 12290
rect 11167 11456 11487 12054
rect 11167 11392 11175 11456
rect 11239 11392 11255 11456
rect 11319 11392 11335 11456
rect 11399 11392 11415 11456
rect 11479 11392 11487 11456
rect 11167 10368 11487 11392
rect 11167 10304 11175 10368
rect 11239 10304 11255 10368
rect 11319 10304 11335 10368
rect 11399 10304 11415 10368
rect 11479 10304 11487 10368
rect 11167 9434 11487 10304
rect 11167 9280 11209 9434
rect 11445 9280 11487 9434
rect 11167 9216 11175 9280
rect 11479 9216 11487 9280
rect 11167 9198 11209 9216
rect 11445 9198 11487 9216
rect 11167 8192 11487 9198
rect 11167 8128 11175 8192
rect 11239 8128 11255 8192
rect 11319 8128 11335 8192
rect 11399 8128 11415 8192
rect 11479 8128 11487 8192
rect 11167 7104 11487 8128
rect 11167 7040 11175 7104
rect 11239 7040 11255 7104
rect 11319 7040 11335 7104
rect 11399 7040 11415 7104
rect 11479 7040 11487 7104
rect 11167 6578 11487 7040
rect 11167 6342 11209 6578
rect 11445 6342 11487 6578
rect 11167 6016 11487 6342
rect 11167 5952 11175 6016
rect 11239 5952 11255 6016
rect 11319 5952 11335 6016
rect 11399 5952 11415 6016
rect 11479 5952 11487 6016
rect 11167 4928 11487 5952
rect 11167 4864 11175 4928
rect 11239 4864 11255 4928
rect 11319 4864 11335 4928
rect 11399 4864 11415 4928
rect 11479 4864 11487 4928
rect 11167 3840 11487 4864
rect 11167 3776 11175 3840
rect 11239 3776 11255 3840
rect 11319 3776 11335 3840
rect 11399 3776 11415 3840
rect 11479 3776 11487 3840
rect 11167 3722 11487 3776
rect 11167 3486 11209 3722
rect 11445 3486 11487 3722
rect 11167 2752 11487 3486
rect 11167 2688 11175 2752
rect 11239 2688 11255 2752
rect 11319 2688 11335 2752
rect 11399 2688 11415 2752
rect 11479 2688 11487 2752
rect 11167 2128 11487 2688
rect 11827 13088 12147 13648
rect 11827 13024 11835 13088
rect 11899 13024 11915 13088
rect 11979 13024 11995 13088
rect 12059 13024 12075 13088
rect 12139 13024 12147 13088
rect 11827 12950 12147 13024
rect 11827 12714 11869 12950
rect 12105 12714 12147 12950
rect 11827 12000 12147 12714
rect 11827 11936 11835 12000
rect 11899 11936 11915 12000
rect 11979 11936 11995 12000
rect 12059 11936 12075 12000
rect 12139 11936 12147 12000
rect 11827 10912 12147 11936
rect 11827 10848 11835 10912
rect 11899 10848 11915 10912
rect 11979 10848 11995 10912
rect 12059 10848 12075 10912
rect 12139 10848 12147 10912
rect 11827 10094 12147 10848
rect 11827 9858 11869 10094
rect 12105 9858 12147 10094
rect 11827 9824 12147 9858
rect 11827 9760 11835 9824
rect 11899 9760 11915 9824
rect 11979 9760 11995 9824
rect 12059 9760 12075 9824
rect 12139 9760 12147 9824
rect 11827 8736 12147 9760
rect 11827 8672 11835 8736
rect 11899 8672 11915 8736
rect 11979 8672 11995 8736
rect 12059 8672 12075 8736
rect 12139 8672 12147 8736
rect 11827 7648 12147 8672
rect 11827 7584 11835 7648
rect 11899 7584 11915 7648
rect 11979 7584 11995 7648
rect 12059 7584 12075 7648
rect 12139 7584 12147 7648
rect 11827 7238 12147 7584
rect 11827 7002 11869 7238
rect 12105 7002 12147 7238
rect 11827 6560 12147 7002
rect 11827 6496 11835 6560
rect 11899 6496 11915 6560
rect 11979 6496 11995 6560
rect 12059 6496 12075 6560
rect 12139 6496 12147 6560
rect 11827 5472 12147 6496
rect 11827 5408 11835 5472
rect 11899 5408 11915 5472
rect 11979 5408 11995 5472
rect 12059 5408 12075 5472
rect 12139 5408 12147 5472
rect 11827 4384 12147 5408
rect 11827 4320 11835 4384
rect 11899 4382 11915 4384
rect 11979 4382 11995 4384
rect 12059 4382 12075 4384
rect 12139 4320 12147 4384
rect 11827 4146 11869 4320
rect 12105 4146 12147 4320
rect 11827 3296 12147 4146
rect 11827 3232 11835 3296
rect 11899 3232 11915 3296
rect 11979 3232 11995 3296
rect 12059 3232 12075 3296
rect 12139 3232 12147 3296
rect 11827 2208 12147 3232
rect 11827 2144 11835 2208
rect 11899 2144 11915 2208
rect 11979 2144 11995 2208
rect 12059 2144 12075 2208
rect 12139 2144 12147 2208
rect 11827 2128 12147 2144
<< via4 >>
rect 2446 12054 2682 12290
rect 2446 9280 2682 9434
rect 2446 9216 2476 9280
rect 2476 9216 2492 9280
rect 2492 9216 2556 9280
rect 2556 9216 2572 9280
rect 2572 9216 2636 9280
rect 2636 9216 2652 9280
rect 2652 9216 2682 9280
rect 2446 9198 2682 9216
rect 2446 6342 2682 6578
rect 2446 3486 2682 3722
rect 3106 12714 3342 12950
rect 3106 9858 3342 10094
rect 3106 7002 3342 7238
rect 3106 4320 3136 4382
rect 3136 4320 3152 4382
rect 3152 4320 3216 4382
rect 3216 4320 3232 4382
rect 3232 4320 3296 4382
rect 3296 4320 3312 4382
rect 3312 4320 3342 4382
rect 3106 4146 3342 4320
rect 5367 12054 5603 12290
rect 5367 9280 5603 9434
rect 5367 9216 5397 9280
rect 5397 9216 5413 9280
rect 5413 9216 5477 9280
rect 5477 9216 5493 9280
rect 5493 9216 5557 9280
rect 5557 9216 5573 9280
rect 5573 9216 5603 9280
rect 5367 9198 5603 9216
rect 5367 6342 5603 6578
rect 5367 3486 5603 3722
rect 6027 12714 6263 12950
rect 6027 9858 6263 10094
rect 6027 7002 6263 7238
rect 6027 4320 6057 4382
rect 6057 4320 6073 4382
rect 6073 4320 6137 4382
rect 6137 4320 6153 4382
rect 6153 4320 6217 4382
rect 6217 4320 6233 4382
rect 6233 4320 6263 4382
rect 6027 4146 6263 4320
rect 8288 12054 8524 12290
rect 8288 9280 8524 9434
rect 8288 9216 8318 9280
rect 8318 9216 8334 9280
rect 8334 9216 8398 9280
rect 8398 9216 8414 9280
rect 8414 9216 8478 9280
rect 8478 9216 8494 9280
rect 8494 9216 8524 9280
rect 8288 9198 8524 9216
rect 8288 6342 8524 6578
rect 8288 3486 8524 3722
rect 8948 12714 9184 12950
rect 8948 9858 9184 10094
rect 8948 7002 9184 7238
rect 8948 4320 8978 4382
rect 8978 4320 8994 4382
rect 8994 4320 9058 4382
rect 9058 4320 9074 4382
rect 9074 4320 9138 4382
rect 9138 4320 9154 4382
rect 9154 4320 9184 4382
rect 8948 4146 9184 4320
rect 11209 12054 11445 12290
rect 11209 9280 11445 9434
rect 11209 9216 11239 9280
rect 11239 9216 11255 9280
rect 11255 9216 11319 9280
rect 11319 9216 11335 9280
rect 11335 9216 11399 9280
rect 11399 9216 11415 9280
rect 11415 9216 11445 9280
rect 11209 9198 11445 9216
rect 11209 6342 11445 6578
rect 11209 3486 11445 3722
rect 11869 12714 12105 12950
rect 11869 9858 12105 10094
rect 11869 7002 12105 7238
rect 11869 4320 11899 4382
rect 11899 4320 11915 4382
rect 11915 4320 11979 4382
rect 11979 4320 11995 4382
rect 11995 4320 12059 4382
rect 12059 4320 12075 4382
rect 12075 4320 12105 4382
rect 11869 4146 12105 4320
<< metal5 >>
rect 1056 12950 12836 12992
rect 1056 12714 3106 12950
rect 3342 12714 6027 12950
rect 6263 12714 8948 12950
rect 9184 12714 11869 12950
rect 12105 12714 12836 12950
rect 1056 12672 12836 12714
rect 1056 12290 12836 12332
rect 1056 12054 2446 12290
rect 2682 12054 5367 12290
rect 5603 12054 8288 12290
rect 8524 12054 11209 12290
rect 11445 12054 12836 12290
rect 1056 12012 12836 12054
rect 1056 10094 12836 10136
rect 1056 9858 3106 10094
rect 3342 9858 6027 10094
rect 6263 9858 8948 10094
rect 9184 9858 11869 10094
rect 12105 9858 12836 10094
rect 1056 9816 12836 9858
rect 1056 9434 12836 9476
rect 1056 9198 2446 9434
rect 2682 9198 5367 9434
rect 5603 9198 8288 9434
rect 8524 9198 11209 9434
rect 11445 9198 12836 9434
rect 1056 9156 12836 9198
rect 1056 7238 12836 7280
rect 1056 7002 3106 7238
rect 3342 7002 6027 7238
rect 6263 7002 8948 7238
rect 9184 7002 11869 7238
rect 12105 7002 12836 7238
rect 1056 6960 12836 7002
rect 1056 6578 12836 6620
rect 1056 6342 2446 6578
rect 2682 6342 5367 6578
rect 5603 6342 8288 6578
rect 8524 6342 11209 6578
rect 11445 6342 12836 6578
rect 1056 6300 12836 6342
rect 1056 4382 12836 4424
rect 1056 4146 3106 4382
rect 3342 4146 6027 4382
rect 6263 4146 8948 4382
rect 9184 4146 11869 4382
rect 12105 4146 12836 4382
rect 1056 4104 12836 4146
rect 1056 3722 12836 3764
rect 1056 3486 2446 3722
rect 2682 3486 5367 3722
rect 5603 3486 8288 3722
rect 8524 3486 11209 3722
rect 11445 3486 12836 3722
rect 1056 3444 12836 3486
use sky130_fd_sc_hd__inv_2  _114_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _115_
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _116_
timestamp 1688980957
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _117_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 2300 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _118_
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _119_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4048 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _120_
timestamp 1688980957
transform 1 0 4416 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _121_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 5336 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _122_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _123_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8648 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _124_
timestamp 1688980957
transform -1 0 8188 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _125_
timestamp 1688980957
transform -1 0 6624 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _126_
timestamp 1688980957
transform -1 0 5888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_4  _127_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7268 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__nor3_1  _128_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7544 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _129_
timestamp 1688980957
transform -1 0 8096 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _130_
timestamp 1688980957
transform -1 0 10120 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_2  _131_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7636 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _132_
timestamp 1688980957
transform -1 0 2024 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _133_
timestamp 1688980957
transform -1 0 4140 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _134_
timestamp 1688980957
transform -1 0 4600 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_2  _135_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4324 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _136_
timestamp 1688980957
transform -1 0 3588 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _137_
timestamp 1688980957
transform -1 0 4876 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _138_
timestamp 1688980957
transform -1 0 6256 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_2  _139_
timestamp 1688980957
transform 1 0 3956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor4_2  _140_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7820 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _141_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9384 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _142_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11040 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _143_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2116 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _144_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _145_
timestamp 1688980957
transform -1 0 5704 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _146_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 2208 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _147_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3680 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _148_
timestamp 1688980957
transform 1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _149_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _150_
timestamp 1688980957
transform -1 0 1840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_1  _151_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2576 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _152_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8464 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _153_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9016 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _154_
timestamp 1688980957
transform -1 0 9016 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _155_
timestamp 1688980957
transform -1 0 10488 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _156_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6808 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_2  _157_
timestamp 1688980957
transform 1 0 7636 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_4  _158_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6532 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__nand4_4  _159_
timestamp 1688980957
transform -1 0 8832 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_1  _160_
timestamp 1688980957
transform -1 0 7452 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _161_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5336 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _162_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3864 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_2  _163_
timestamp 1688980957
transform 1 0 5612 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _164_
timestamp 1688980957
transform -1 0 6256 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _165_
timestamp 1688980957
transform 1 0 5060 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _166_
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _167_
timestamp 1688980957
transform 1 0 2024 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _168_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4508 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _169_
timestamp 1688980957
transform 1 0 4968 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _170_
timestamp 1688980957
transform -1 0 7820 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _171_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7728 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _172_
timestamp 1688980957
transform -1 0 8832 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _173_
timestamp 1688980957
transform 1 0 5244 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _174_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 6256 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _175_
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2ai_2  _176_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7912 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_1  _177_
timestamp 1688980957
transform -1 0 5060 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_1  _178_
timestamp 1688980957
transform -1 0 6808 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a22oi_2  _179_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6072 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _180_
timestamp 1688980957
transform 1 0 5612 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o22ai_1  _181_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7084 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _182_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9476 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _183_
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _184_
timestamp 1688980957
transform -1 0 9200 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2ai_1  _185_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8740 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_1  _186_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4232 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _187_
timestamp 1688980957
transform -1 0 3956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _188_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4692 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _189_
timestamp 1688980957
transform 1 0 5612 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _190_
timestamp 1688980957
transform 1 0 10212 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _191_
timestamp 1688980957
transform 1 0 3496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor4_1  _192_
timestamp 1688980957
transform -1 0 8648 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o22ai_1  _193_
timestamp 1688980957
transform 1 0 9568 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _194_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8832 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _195_
timestamp 1688980957
transform -1 0 10488 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _197_
timestamp 1688980957
transform 1 0 5336 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _198_
timestamp 1688980957
transform -1 0 6256 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _199_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7820 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _200_
timestamp 1688980957
transform -1 0 10028 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _201_
timestamp 1688980957
transform 1 0 10948 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _202_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9016 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _203_
timestamp 1688980957
transform -1 0 3036 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _204_
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _205_
timestamp 1688980957
transform -1 0 2852 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _206_
timestamp 1688980957
transform -1 0 5244 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _207_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _208_
timestamp 1688980957
transform -1 0 5980 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _209_
timestamp 1688980957
transform 1 0 6716 0 1 2176
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _210_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7820 0 -1 3264
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _211_
timestamp 1688980957
transform 1 0 9200 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _212_
timestamp 1688980957
transform -1 0 8556 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _213__31 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3036 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _213_
timestamp 1688980957
transform 1 0 4416 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _214__30
timestamp 1688980957
transform 1 0 4324 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _214_
timestamp 1688980957
transform 1 0 4324 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _215__29
timestamp 1688980957
transform -1 0 5152 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _215_
timestamp 1688980957
transform 1 0 4600 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _216__28
timestamp 1688980957
transform -1 0 2392 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _216_
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _217__27
timestamp 1688980957
transform -1 0 6164 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _217_
timestamp 1688980957
transform 1 0 4968 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _218__26
timestamp 1688980957
transform 1 0 4508 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _218_
timestamp 1688980957
transform 1 0 4784 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _219__25
timestamp 1688980957
transform 1 0 2024 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _219_
timestamp 1688980957
transform 1 0 2024 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _220__24
timestamp 1688980957
transform 1 0 6624 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _220_
timestamp 1688980957
transform 1 0 6900 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _221__23
timestamp 1688980957
transform 1 0 2300 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _221_
timestamp 1688980957
transform 1 0 2208 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _222__22
timestamp 1688980957
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _222_
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _223__21
timestamp 1688980957
transform 1 0 6900 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _223_
timestamp 1688980957
transform 1 0 7176 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _224__20
timestamp 1688980957
transform -1 0 6716 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _224_
timestamp 1688980957
transform 1 0 5796 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _225__19
timestamp 1688980957
transform -1 0 3036 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _225_
timestamp 1688980957
transform 1 0 2208 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _226_
timestamp 1688980957
transform 1 0 6440 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _226__18
timestamp 1688980957
transform -1 0 6992 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _227__17
timestamp 1688980957
transform -1 0 3772 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _227_
timestamp 1688980957
transform 1 0 3312 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _228_
timestamp 1688980957
transform 1 0 3772 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _228__16
timestamp 1688980957
transform -1 0 4324 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _229__15
timestamp 1688980957
transform -1 0 9200 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _229_
timestamp 1688980957
transform 1 0 8372 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _230__14
timestamp 1688980957
transform 1 0 4876 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _230_
timestamp 1688980957
transform 1 0 4784 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _231__13
timestamp 1688980957
transform -1 0 9476 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _231_
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _232__12
timestamp 1688980957
transform -1 0 7452 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _232_
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _233__11
timestamp 1688980957
transform -1 0 2116 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _233_
timestamp 1688980957
transform 1 0 1564 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _234__10
timestamp 1688980957
transform -1 0 7176 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _234_
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _235__9
timestamp 1688980957
transform 1 0 1472 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _235_
timestamp 1688980957
transform 1 0 2208 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _236__8
timestamp 1688980957
transform -1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _236_
timestamp 1688980957
transform 1 0 5428 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _237__7
timestamp 1688980957
transform 1 0 1748 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _237_
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _238__6
timestamp 1688980957
transform -1 0 7176 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _238_
timestamp 1688980957
transform 1 0 6624 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _239__5
timestamp 1688980957
transform -1 0 6624 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _239_
timestamp 1688980957
transform 1 0 5152 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _240_
timestamp 1688980957
transform 1 0 4416 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _241_
timestamp 1688980957
transform 1 0 8740 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5796 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1688980957
transform -1 0 4416 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1688980957
transform 1 0 5244 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1688980957
transform -1 0 4416 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1688980957
transform 1 0 5244 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1932 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_50 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5704 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_54
timestamp 1688980957
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_60
timestamp 1688980957
transform 1 0 6624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_78
timestamp 1688980957
transform 1 0 8280 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_88 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9200 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_100
timestamp 1688980957
transform 1 0 10304 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_113 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_65
timestamp 1688980957
transform 1 0 7084 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_92
timestamp 1688980957
transform 1 0 9568 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_104
timestamp 1688980957
transform 1 0 10672 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_121 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12236 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_43
timestamp 1688980957
transform 1 0 5060 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_73
timestamp 1688980957
transform 1 0 7820 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_82
timestamp 1688980957
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_91
timestamp 1688980957
transform 1 0 9476 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_102
timestamp 1688980957
transform 1 0 10488 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_114
timestamp 1688980957
transform 1 0 11592 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_122
timestamp 1688980957
transform 1 0 12328 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_74
timestamp 1688980957
transform 1 0 7912 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_121
timestamp 1688980957
transform 1 0 12236 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_19
timestamp 1688980957
transform 1 0 2852 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_64
timestamp 1688980957
transform 1 0 6992 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_100
timestamp 1688980957
transform 1 0 10304 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_112
timestamp 1688980957
transform 1 0 11408 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_9
timestamp 1688980957
transform 1 0 1932 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_86 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9016 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_102
timestamp 1688980957
transform 1 0 10488 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_110
timestamp 1688980957
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_121
timestamp 1688980957
transform 1 0 12236 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_82
timestamp 1688980957
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_113
timestamp 1688980957
transform 1 0 11500 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_73
timestamp 1688980957
transform 1 0 7820 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_121
timestamp 1688980957
transform 1 0 12236 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_10
timestamp 1688980957
transform 1 0 2024 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_34
timestamp 1688980957
transform 1 0 4232 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_9
timestamp 1688980957
transform 1 0 1932 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_52
timestamp 1688980957
transform 1 0 5888 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_110
timestamp 1688980957
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_121
timestamp 1688980957
transform 1 0 12236 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_19
timestamp 1688980957
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_33
timestamp 1688980957
transform 1 0 4140 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_38
timestamp 1688980957
transform 1 0 4600 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_42
timestamp 1688980957
transform 1 0 4968 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_80
timestamp 1688980957
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_101
timestamp 1688980957
transform 1 0 10396 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_113
timestamp 1688980957
transform 1 0 11500 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_76
timestamp 1688980957
transform 1 0 8096 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_98
timestamp 1688980957
transform 1 0 10120 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_110
timestamp 1688980957
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_121
timestamp 1688980957
transform 1 0 12236 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_7
timestamp 1688980957
transform 1 0 1748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_14
timestamp 1688980957
transform 1 0 2392 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_22
timestamp 1688980957
transform 1 0 3128 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_45
timestamp 1688980957
transform 1 0 5244 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_69
timestamp 1688980957
transform 1 0 7452 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_79
timestamp 1688980957
transform 1 0 8372 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_91
timestamp 1688980957
transform 1 0 9476 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_103
timestamp 1688980957
transform 1 0 10580 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_115
timestamp 1688980957
transform 1 0 11684 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_123
timestamp 1688980957
transform 1 0 12420 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_21
timestamp 1688980957
transform 1 0 3036 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_60
timestamp 1688980957
transform 1 0 6624 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_70
timestamp 1688980957
transform 1 0 7544 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_82
timestamp 1688980957
transform 1 0 8648 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_94
timestamp 1688980957
transform 1 0 9752 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_106
timestamp 1688980957
transform 1 0 10856 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_121
timestamp 1688980957
transform 1 0 12236 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_11
timestamp 1688980957
transform 1 0 2116 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_35
timestamp 1688980957
transform 1 0 4324 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_76
timestamp 1688980957
transform 1 0 8096 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1688980957
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1688980957
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_121
timestamp 1688980957
transform 1 0 12236 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_15
timestamp 1688980957
transform 1 0 2484 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_23
timestamp 1688980957
transform 1 0 3220 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_45
timestamp 1688980957
transform 1 0 5244 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_49
timestamp 1688980957
transform 1 0 5612 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_53
timestamp 1688980957
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1688980957
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1688980957
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1688980957
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1688980957
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1688980957
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_121
timestamp 1688980957
transform 1 0 12236 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1688980957
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_41
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_58
timestamp 1688980957
transform 1 0 6440 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_62
timestamp 1688980957
transform 1 0 6808 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_79
timestamp 1688980957
transform 1 0 8372 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1688980957
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1688980957
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 1688980957
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_121
timestamp 1688980957
transform 1 0 12236 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1688980957
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_27
timestamp 1688980957
transform 1 0 3588 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_35
timestamp 1688980957
transform 1 0 4324 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_85
timestamp 1688980957
transform 1 0 8924 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_97
timestamp 1688980957
transform 1 0 10028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_109
timestamp 1688980957
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_121
timestamp 1688980957
transform 1 0 12236 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1688980957
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1688980957
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 1688980957
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_121
timestamp 1688980957
transform 1 0 12236 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1688980957
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_27
timestamp 1688980957
transform 1 0 3588 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_54
timestamp 1688980957
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_77
timestamp 1688980957
transform 1 0 8188 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_89
timestamp 1688980957
transform 1 0 9292 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_101
timestamp 1688980957
transform 1 0 10396 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_109
timestamp 1688980957
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_121
timestamp 1688980957
transform 1 0 12236 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1688980957
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_44
timestamp 1688980957
transform 1 0 5152 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_48
timestamp 1688980957
transform 1 0 5520 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_55
timestamp 1688980957
transform 1 0 6164 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_57
timestamp 1688980957
transform 1 0 6348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_64
timestamp 1688980957
transform 1 0 6992 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_76
timestamp 1688980957
transform 1 0 8096 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1688980957
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_109
timestamp 1688980957
transform 1 0 11132 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_113
timestamp 1688980957
transform 1 0 11500 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4508 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform -1 0 3680 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform 1 0 2300 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform -1 0 3588 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform -1 0 7820 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform -1 0 8648 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform -1 0 3772 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform 1 0 3772 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform -1 0 11224 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform 1 0 9476 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform -1 0 5796 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform -1 0 10948 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1688980957
transform 1 0 12236 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1688980957
transform 1 0 12236 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  max_cap4 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 11500 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 1932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 12788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 12788 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 12788 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 12788 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 12788 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 12788 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 12788 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 12788 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 12788 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 12788 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 12788 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 12788 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 12788 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 12788 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 12788 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 12788 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 12788 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 12788 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 12788 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 12788 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 12788 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 6256 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 11408 0 1 13056
box -38 -48 130 592
<< labels >>
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 PWM_OUT
port 0 nsew signal tristate
flabel metal4 s 3064 2128 3384 13648 0 FreeSans 1920 90 0 0 VGND
port 1 nsew ground bidirectional
flabel metal4 s 5985 2128 6305 13648 0 FreeSans 1920 90 0 0 VGND
port 1 nsew ground bidirectional
flabel metal4 s 8906 2128 9226 13648 0 FreeSans 1920 90 0 0 VGND
port 1 nsew ground bidirectional
flabel metal4 s 11827 2128 12147 13648 0 FreeSans 1920 90 0 0 VGND
port 1 nsew ground bidirectional
flabel metal5 s 1056 4104 12836 4424 0 FreeSans 2560 0 0 0 VGND
port 1 nsew ground bidirectional
flabel metal5 s 1056 6960 12836 7280 0 FreeSans 2560 0 0 0 VGND
port 1 nsew ground bidirectional
flabel metal5 s 1056 9816 12836 10136 0 FreeSans 2560 0 0 0 VGND
port 1 nsew ground bidirectional
flabel metal5 s 1056 12672 12836 12992 0 FreeSans 2560 0 0 0 VGND
port 1 nsew ground bidirectional
flabel metal4 s 2404 2128 2724 13648 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal4 s 5325 2128 5645 13648 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal4 s 8246 2128 8566 13648 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal4 s 11167 2128 11487 13648 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal5 s 1056 3444 12836 3764 0 FreeSans 2560 0 0 0 VPWR
port 2 nsew power bidirectional
flabel metal5 s 1056 6300 12836 6620 0 FreeSans 2560 0 0 0 VPWR
port 2 nsew power bidirectional
flabel metal5 s 1056 9156 12836 9476 0 FreeSans 2560 0 0 0 VPWR
port 2 nsew power bidirectional
flabel metal5 s 1056 12012 12836 12332 0 FreeSans 2560 0 0 0 VPWR
port 2 nsew power bidirectional
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 clk
port 3 nsew signal input
flabel metal2 s 13542 15266 13598 16066 0 FreeSans 224 90 0 0 decrease_duty
port 4 nsew signal input
flabel metal3 s 13122 688 13922 808 0 FreeSans 480 0 0 0 increase_duty
port 5 nsew signal input
rlabel metal1 6946 13056 6946 13056 0 VGND
rlabel metal1 6946 13600 6946 13600 0 VPWR
rlabel metal1 4462 4148 4462 4148 0 DUTY_CYCLE\[0\]
rlabel metal2 8970 4879 8970 4879 0 DUTY_CYCLE\[1\]
rlabel metal2 4738 4930 4738 4930 0 DUTY_CYCLE\[2\]
rlabel metal2 8418 5423 8418 5423 0 DUTY_CYCLE\[3\]
rlabel metal1 10350 3434 10350 3434 0 PWM_DFF1.Q
rlabel metal1 5796 6154 5796 6154 0 PWM_DFF2.Q
rlabel metal1 9200 5134 9200 5134 0 PWM_DFF3.Q
rlabel metal2 10442 5593 10442 5593 0 PWM_DFF4.Q
rlabel metal2 46 1554 46 1554 0 PWM_OUT
rlabel metal1 9747 5678 9747 5678 0 _000_
rlabel metal2 3726 4284 3726 4284 0 _001_
rlabel via1 1697 4522 1697 4522 0 _002_
rlabel metal1 2806 2924 2806 2924 0 _003_
rlabel metal1 2852 2618 2852 2618 0 _004_
rlabel metal1 6210 2958 6210 2958 0 _005_
rlabel metal1 5060 4658 5060 4658 0 _006_
rlabel via1 7028 2414 7028 2414 0 _007_
rlabel metal1 8372 2958 8372 2958 0 _008_
rlabel metal1 9793 4114 9793 4114 0 _009_
rlabel metal1 7778 6766 7778 6766 0 _010_
rlabel metal2 7130 7174 7130 7174 0 _038_
rlabel metal1 10023 7446 10023 7446 0 _039_
rlabel metal2 9982 8738 9982 8738 0 _040_
rlabel metal1 7820 7854 7820 7854 0 _041_
rlabel metal1 2323 6426 2323 6426 0 _042_
rlabel metal2 4646 7276 4646 7276 0 _043_
rlabel metal2 4370 7242 4370 7242 0 _044_
rlabel metal1 5382 5644 5382 5644 0 _045_
rlabel metal2 4002 8262 4002 8262 0 _046_
rlabel metal1 4922 8602 4922 8602 0 _047_
rlabel metal1 4646 8364 4646 8364 0 _048_
rlabel metal1 5110 5678 5110 5678 0 _049_
rlabel metal1 9338 6902 9338 6902 0 _050_
rlabel metal1 9476 5338 9476 5338 0 _051_
rlabel metal1 3312 2278 3312 2278 0 _052_
rlabel metal1 4692 2278 4692 2278 0 _053_
rlabel metal1 3220 4182 3220 4182 0 _054_
rlabel metal1 2162 5032 2162 5032 0 _055_
rlabel metal1 2484 2482 2484 2482 0 _056_
rlabel metal1 7921 5678 7921 5678 0 _057_
rlabel metal2 7866 5984 7866 5984 0 _058_
rlabel metal1 7912 5066 7912 5066 0 _059_
rlabel metal1 7314 5236 7314 5236 0 _060_
rlabel metal1 7682 5168 7682 5168 0 _061_
rlabel metal1 5842 4114 5842 4114 0 _062_
rlabel metal1 10994 6222 10994 6222 0 _063_
rlabel metal1 9246 2414 9246 2414 0 _064_
rlabel metal1 5750 2958 5750 2958 0 _065_
rlabel metal1 5658 5712 5658 5712 0 _066_
rlabel metal1 6026 5270 6026 5270 0 _067_
rlabel metal1 5244 4114 5244 4114 0 _068_
rlabel metal1 5198 4250 5198 4250 0 _069_
rlabel metal1 2392 5202 2392 5202 0 _070_
rlabel metal2 2070 4896 2070 4896 0 _071_
rlabel metal1 5474 4692 5474 4692 0 _072_
rlabel metal2 6670 3519 6670 3519 0 _073_
rlabel metal1 8096 5882 8096 5882 0 _074_
rlabel metal1 8326 5644 8326 5644 0 _075_
rlabel metal1 5704 5882 5704 5882 0 _076_
rlabel viali 8689 6222 8689 6222 0 _077_
rlabel metal1 8786 6324 8786 6324 0 _078_
rlabel metal1 8234 4148 8234 4148 0 _079_
rlabel metal1 7038 2856 7038 2856 0 _080_
rlabel metal1 6578 4624 6578 4624 0 _081_
rlabel metal1 6670 4522 6670 4522 0 _082_
rlabel metal1 6854 3026 6854 3026 0 _083_
rlabel metal1 8786 2380 8786 2380 0 _084_
rlabel metal2 8694 4284 8694 4284 0 _085_
rlabel metal1 8602 4080 8602 4080 0 _086_
rlabel metal1 8510 3910 8510 3910 0 _087_
rlabel metal1 4416 6630 4416 6630 0 _088_
rlabel metal1 3910 8364 3910 8364 0 _089_
rlabel metal2 3542 6528 3542 6528 0 _090_
rlabel metal1 7682 6290 7682 6290 0 _091_
rlabel metal1 10028 4590 10028 4590 0 _092_
rlabel metal1 7033 6222 7033 6222 0 _093_
rlabel metal2 9890 5168 9890 5168 0 _094_
rlabel metal1 9154 2278 9154 2278 0 _095_
rlabel metal1 10350 3706 10350 3706 0 _096_
rlabel metal1 5980 7378 5980 7378 0 _097_
rlabel metal1 10534 6630 10534 6630 0 _098_
rlabel metal1 5658 2278 5658 2278 0 _099_
rlabel viali 4738 3027 4738 3027 0 _100_
rlabel metal1 2438 3026 2438 3026 0 _101_
rlabel via1 4554 3179 4554 3179 0 _102_
rlabel metal1 6532 3162 6532 3162 0 _103_
rlabel metal1 4554 3502 4554 3502 0 _104_
rlabel metal1 5290 3060 5290 3060 0 _105_
rlabel metal1 3358 2516 3358 2516 0 _106_
rlabel metal1 8740 11866 8740 11866 0 _107_
rlabel metal2 8142 12410 8142 12410 0 _108_
rlabel metal1 7084 11866 7084 11866 0 _109_
rlabel metal1 6532 13362 6532 13362 0 _110_
rlabel metal2 8142 8925 8142 8925 0 _111_
rlabel metal1 7590 8942 7590 8942 0 _112_
rlabel metal2 7958 8772 7958 8772 0 _113_
rlabel metal2 4094 14433 4094 14433 0 clk
rlabel metal1 4876 7446 4876 7446 0 clknet_0_clk
rlabel metal1 2070 6154 2070 6154 0 clknet_2_0__leaf_clk
rlabel metal1 5980 2482 5980 2482 0 clknet_2_1__leaf_clk
rlabel metal1 1518 8398 1518 8398 0 clknet_2_2__leaf_clk
rlabel metal1 8418 8330 8418 8330 0 clknet_2_3__leaf_clk
rlabel metal2 2254 3196 2254 3196 0 counter_PWM\[0\]
rlabel metal1 2484 4454 2484 4454 0 counter_PWM\[1\]
rlabel metal1 2530 2958 2530 2958 0 counter_PWM\[2\]
rlabel metal2 3818 2176 3818 2176 0 counter_PWM\[3\]
rlabel metal1 5198 6834 5198 6834 0 counter_debounce\[0\]
rlabel metal1 4508 8806 4508 8806 0 counter_debounce\[10\]
rlabel metal1 8648 11730 8648 11730 0 counter_debounce\[11\]
rlabel metal1 7590 12410 7590 12410 0 counter_debounce\[12\]
rlabel metal1 4094 9962 4094 9962 0 counter_debounce\[13\]
rlabel metal1 8142 12784 8142 12784 0 counter_debounce\[14\]
rlabel metal2 4738 9860 4738 9860 0 counter_debounce\[15\]
rlabel metal1 4830 10064 4830 10064 0 counter_debounce\[16\]
rlabel metal1 9844 8466 9844 8466 0 counter_debounce\[17\]
rlabel metal1 6210 8534 6210 8534 0 counter_debounce\[18\]
rlabel metal1 10212 8058 10212 8058 0 counter_debounce\[19\]
rlabel metal1 4692 7854 4692 7854 0 counter_debounce\[1\]
rlabel metal1 7820 7514 7820 7514 0 counter_debounce\[20\]
rlabel metal1 3542 8432 3542 8432 0 counter_debounce\[21\]
rlabel metal1 8050 8500 8050 8500 0 counter_debounce\[22\]
rlabel metal1 1794 6324 1794 6324 0 counter_debounce\[23\]
rlabel metal1 7038 9146 7038 9146 0 counter_debounce\[24\]
rlabel metal1 1978 6188 1978 6188 0 counter_debounce\[25\]
rlabel metal1 7774 9554 7774 9554 0 counter_debounce\[26\]
rlabel metal2 7406 9724 7406 9724 0 counter_debounce\[27\]
rlabel metal2 5704 12852 5704 12852 0 counter_debounce\[2\]
rlabel metal1 5980 12954 5980 12954 0 counter_debounce\[3\]
rlabel metal1 3082 8058 3082 8058 0 counter_debounce\[4\]
rlabel metal2 6394 11526 6394 11526 0 counter_debounce\[5\]
rlabel metal1 6578 11696 6578 11696 0 counter_debounce\[6\]
rlabel metal1 3864 6834 3864 6834 0 counter_debounce\[7\]
rlabel metal1 8602 11322 8602 11322 0 counter_debounce\[8\]
rlabel metal1 4002 6970 4002 6970 0 counter_debounce\[9\]
rlabel metal1 12466 13328 12466 13328 0 decrease_duty
rlabel metal1 12650 2414 12650 2414 0 increase_duty
rlabel metal1 10902 6834 10902 6834 0 net1
rlabel metal1 6803 8534 6803 8534 0 net10
rlabel via1 1881 8534 1881 8534 0 net11
rlabel metal1 6941 7446 6941 7446 0 net12
rlabel metal1 9287 7786 9287 7786 0 net13
rlabel via1 5101 9622 5101 9622 0 net14
rlabel metal1 8735 8534 8735 8534 0 net15
rlabel metal2 4094 10438 4094 10438 0 net16
rlabel via1 3629 9554 3629 9554 0 net17
rlabel via1 6757 12818 6757 12818 0 net18
rlabel metal2 2806 9724 2806 9724 0 net19
rlabel metal1 11132 3502 11132 3502 0 net2
rlabel metal2 6440 12852 6440 12852 0 net20
rlabel metal1 7304 11730 7304 11730 0 net21
rlabel metal1 3854 8942 3854 8942 0 net22
rlabel metal1 2422 6698 2422 6698 0 net23
rlabel metal1 7120 11118 7120 11118 0 net24
rlabel metal2 2300 6596 2300 6596 0 net25
rlabel metal1 4825 11662 4825 11662 0 net26
rlabel metal1 6256 13430 6256 13430 0 net27
rlabel metal1 1927 7854 1927 7854 0 net28
rlabel via1 4917 12886 4917 12886 0 net29
rlabel metal1 2484 2346 2484 2346 0 net3
rlabel metal2 4554 12517 4554 12517 0 net30
rlabel metal1 4636 7378 4636 7378 0 net31
rlabel metal1 1978 5780 1978 5780 0 net32
rlabel metal1 2672 4182 2672 4182 0 net33
rlabel metal1 6210 2414 6210 2414 0 net34
rlabel metal1 2729 3434 2729 3434 0 net35
rlabel metal1 5566 3060 5566 3060 0 net36
rlabel metal1 7774 3060 7774 3060 0 net37
rlabel metal2 3082 2720 3082 2720 0 net38
rlabel metal1 4696 2414 4696 2414 0 net39
rlabel metal1 11270 5576 11270 5576 0 net4
rlabel metal1 10166 5338 10166 5338 0 net40
rlabel metal1 11270 6324 11270 6324 0 net41
rlabel metal1 7222 6290 7222 6290 0 net42
rlabel metal1 4917 6358 4917 6358 0 net43
rlabel metal2 9614 7072 9614 7072 0 net44
rlabel metal1 6164 9554 6164 9554 0 net5
rlabel metal2 6946 9758 6946 9758 0 net6
rlabel metal1 1978 6698 1978 6698 0 net7
rlabel via1 5745 8874 5745 8874 0 net8
rlabel metal1 2100 5610 2100 5610 0 net9
<< properties >>
string FIXED_BBOX 0 0 13922 16066
<< end >>
